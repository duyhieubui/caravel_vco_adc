// This is the unpowered netlist.
module vco_adc (clk,
    data_valid_out,
    enable_in,
    rst,
    data_out,
    oversample_in,
    phase_in);
 input clk;
 output data_valid_out;
 input enable_in;
 input rst;
 output [31:0] data_out;
 input [9:0] oversample_in;
 input [10:0] phase_in;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net867;
 wire net868;
 wire net87;
 wire net870;
 wire net872;
 wire net873;
 wire net874;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire output_en_reg;
 wire \pr.genblk1[0].pd.ff_reg_0 ;
 wire \pr.genblk1[0].pd.ff_reg_1 ;
 wire \pr.genblk1[10].pd.ff_reg_0 ;
 wire \pr.genblk1[10].pd.ff_reg_1 ;
 wire \pr.genblk1[1].pd.ff_reg_0 ;
 wire \pr.genblk1[1].pd.ff_reg_1 ;
 wire \pr.genblk1[2].pd.ff_reg_0 ;
 wire \pr.genblk1[2].pd.ff_reg_1 ;
 wire \pr.genblk1[3].pd.ff_reg_0 ;
 wire \pr.genblk1[3].pd.ff_reg_1 ;
 wire \pr.genblk1[4].pd.ff_reg_0 ;
 wire \pr.genblk1[4].pd.ff_reg_1 ;
 wire \pr.genblk1[5].pd.ff_reg_0 ;
 wire \pr.genblk1[5].pd.ff_reg_1 ;
 wire \pr.genblk1[6].pd.ff_reg_0 ;
 wire \pr.genblk1[6].pd.ff_reg_1 ;
 wire \pr.genblk1[7].pd.ff_reg_0 ;
 wire \pr.genblk1[7].pd.ff_reg_1 ;
 wire \pr.genblk1[8].pd.ff_reg_0 ;
 wire \pr.genblk1[8].pd.ff_reg_1 ;
 wire \pr.genblk1[9].pd.ff_reg_0 ;
 wire \pr.genblk1[9].pd.ff_reg_1 ;
 wire \scs.acc1[0] ;
 wire \scs.acc1[10] ;
 wire \scs.acc1[11] ;
 wire \scs.acc1[12] ;
 wire \scs.acc1[13] ;
 wire \scs.acc1[14] ;
 wire \scs.acc1[15] ;
 wire \scs.acc1[16] ;
 wire \scs.acc1[17] ;
 wire \scs.acc1[18] ;
 wire \scs.acc1[19] ;
 wire \scs.acc1[1] ;
 wire \scs.acc1[20] ;
 wire \scs.acc1[21] ;
 wire \scs.acc1[22] ;
 wire \scs.acc1[23] ;
 wire \scs.acc1[24] ;
 wire \scs.acc1[25] ;
 wire \scs.acc1[26] ;
 wire \scs.acc1[27] ;
 wire \scs.acc1[28] ;
 wire \scs.acc1[29] ;
 wire \scs.acc1[2] ;
 wire \scs.acc1[30] ;
 wire \scs.acc1[31] ;
 wire \scs.acc1[3] ;
 wire \scs.acc1[4] ;
 wire \scs.acc1[5] ;
 wire \scs.acc1[6] ;
 wire \scs.acc1[7] ;
 wire \scs.acc1[8] ;
 wire \scs.acc1[9] ;
 wire \scs.acc2[0] ;
 wire \scs.acc2[10] ;
 wire \scs.acc2[11] ;
 wire \scs.acc2[12] ;
 wire \scs.acc2[13] ;
 wire \scs.acc2[14] ;
 wire \scs.acc2[15] ;
 wire \scs.acc2[16] ;
 wire \scs.acc2[17] ;
 wire \scs.acc2[18] ;
 wire \scs.acc2[19] ;
 wire \scs.acc2[1] ;
 wire \scs.acc2[20] ;
 wire \scs.acc2[21] ;
 wire \scs.acc2[22] ;
 wire \scs.acc2[23] ;
 wire \scs.acc2[24] ;
 wire \scs.acc2[25] ;
 wire \scs.acc2[26] ;
 wire \scs.acc2[27] ;
 wire \scs.acc2[28] ;
 wire \scs.acc2[29] ;
 wire \scs.acc2[2] ;
 wire \scs.acc2[30] ;
 wire \scs.acc2[31] ;
 wire \scs.acc2[3] ;
 wire \scs.acc2[4] ;
 wire \scs.acc2[5] ;
 wire \scs.acc2[6] ;
 wire \scs.acc2[7] ;
 wire \scs.acc2[8] ;
 wire \scs.acc2[9] ;
 wire \scs.acc3[0] ;
 wire \scs.acc3[10] ;
 wire \scs.acc3[11] ;
 wire \scs.acc3[12] ;
 wire \scs.acc3[13] ;
 wire \scs.acc3[14] ;
 wire \scs.acc3[15] ;
 wire \scs.acc3[16] ;
 wire \scs.acc3[17] ;
 wire \scs.acc3[18] ;
 wire \scs.acc3[19] ;
 wire \scs.acc3[1] ;
 wire \scs.acc3[20] ;
 wire \scs.acc3[21] ;
 wire \scs.acc3[22] ;
 wire \scs.acc3[23] ;
 wire \scs.acc3[24] ;
 wire \scs.acc3[25] ;
 wire \scs.acc3[26] ;
 wire \scs.acc3[27] ;
 wire \scs.acc3[28] ;
 wire \scs.acc3[29] ;
 wire \scs.acc3[2] ;
 wire \scs.acc3[30] ;
 wire \scs.acc3[31] ;
 wire \scs.acc3[3] ;
 wire \scs.acc3[4] ;
 wire \scs.acc3[5] ;
 wire \scs.acc3[6] ;
 wire \scs.acc3[7] ;
 wire \scs.acc3[8] ;
 wire \scs.acc3[9] ;
 wire \scs.acc3_d2[0] ;
 wire \scs.acc3_d2[10] ;
 wire \scs.acc3_d2[11] ;
 wire \scs.acc3_d2[12] ;
 wire \scs.acc3_d2[13] ;
 wire \scs.acc3_d2[14] ;
 wire \scs.acc3_d2[15] ;
 wire \scs.acc3_d2[16] ;
 wire \scs.acc3_d2[17] ;
 wire \scs.acc3_d2[18] ;
 wire \scs.acc3_d2[19] ;
 wire \scs.acc3_d2[1] ;
 wire \scs.acc3_d2[20] ;
 wire \scs.acc3_d2[21] ;
 wire \scs.acc3_d2[22] ;
 wire \scs.acc3_d2[23] ;
 wire \scs.acc3_d2[24] ;
 wire \scs.acc3_d2[25] ;
 wire \scs.acc3_d2[26] ;
 wire \scs.acc3_d2[27] ;
 wire \scs.acc3_d2[28] ;
 wire \scs.acc3_d2[29] ;
 wire \scs.acc3_d2[2] ;
 wire \scs.acc3_d2[30] ;
 wire \scs.acc3_d2[31] ;
 wire \scs.acc3_d2[3] ;
 wire \scs.acc3_d2[4] ;
 wire \scs.acc3_d2[5] ;
 wire \scs.acc3_d2[6] ;
 wire \scs.acc3_d2[7] ;
 wire \scs.acc3_d2[8] ;
 wire \scs.acc3_d2[9] ;
 wire \scs.data_valid_out ;
 wire \scs.decimation_en ;
 wire \scs.diff1[0] ;
 wire \scs.diff1[10] ;
 wire \scs.diff1[11] ;
 wire \scs.diff1[12] ;
 wire \scs.diff1[13] ;
 wire \scs.diff1[14] ;
 wire \scs.diff1[15] ;
 wire \scs.diff1[16] ;
 wire \scs.diff1[17] ;
 wire \scs.diff1[18] ;
 wire \scs.diff1[19] ;
 wire \scs.diff1[1] ;
 wire \scs.diff1[20] ;
 wire \scs.diff1[21] ;
 wire \scs.diff1[22] ;
 wire \scs.diff1[23] ;
 wire \scs.diff1[24] ;
 wire \scs.diff1[25] ;
 wire \scs.diff1[26] ;
 wire \scs.diff1[27] ;
 wire \scs.diff1[28] ;
 wire \scs.diff1[29] ;
 wire \scs.diff1[2] ;
 wire \scs.diff1[30] ;
 wire \scs.diff1[31] ;
 wire \scs.diff1[3] ;
 wire \scs.diff1[4] ;
 wire \scs.diff1[5] ;
 wire \scs.diff1[6] ;
 wire \scs.diff1[7] ;
 wire \scs.diff1[8] ;
 wire \scs.diff1[9] ;
 wire \scs.diff1_d[0] ;
 wire \scs.diff1_d[10] ;
 wire \scs.diff1_d[11] ;
 wire \scs.diff1_d[12] ;
 wire \scs.diff1_d[13] ;
 wire \scs.diff1_d[14] ;
 wire \scs.diff1_d[15] ;
 wire \scs.diff1_d[16] ;
 wire \scs.diff1_d[17] ;
 wire \scs.diff1_d[18] ;
 wire \scs.diff1_d[19] ;
 wire \scs.diff1_d[1] ;
 wire \scs.diff1_d[20] ;
 wire \scs.diff1_d[21] ;
 wire \scs.diff1_d[22] ;
 wire \scs.diff1_d[23] ;
 wire \scs.diff1_d[24] ;
 wire \scs.diff1_d[25] ;
 wire \scs.diff1_d[26] ;
 wire \scs.diff1_d[27] ;
 wire \scs.diff1_d[28] ;
 wire \scs.diff1_d[29] ;
 wire \scs.diff1_d[2] ;
 wire \scs.diff1_d[30] ;
 wire \scs.diff1_d[31] ;
 wire \scs.diff1_d[3] ;
 wire \scs.diff1_d[4] ;
 wire \scs.diff1_d[5] ;
 wire \scs.diff1_d[6] ;
 wire \scs.diff1_d[7] ;
 wire \scs.diff1_d[8] ;
 wire \scs.diff1_d[9] ;
 wire \scs.diff2[0] ;
 wire \scs.diff2[10] ;
 wire \scs.diff2[11] ;
 wire \scs.diff2[12] ;
 wire \scs.diff2[13] ;
 wire \scs.diff2[14] ;
 wire \scs.diff2[15] ;
 wire \scs.diff2[16] ;
 wire \scs.diff2[17] ;
 wire \scs.diff2[18] ;
 wire \scs.diff2[19] ;
 wire \scs.diff2[1] ;
 wire \scs.diff2[20] ;
 wire \scs.diff2[21] ;
 wire \scs.diff2[22] ;
 wire \scs.diff2[23] ;
 wire \scs.diff2[24] ;
 wire \scs.diff2[25] ;
 wire \scs.diff2[26] ;
 wire \scs.diff2[27] ;
 wire \scs.diff2[28] ;
 wire \scs.diff2[29] ;
 wire \scs.diff2[2] ;
 wire \scs.diff2[30] ;
 wire \scs.diff2[31] ;
 wire \scs.diff2[3] ;
 wire \scs.diff2[4] ;
 wire \scs.diff2[5] ;
 wire \scs.diff2[6] ;
 wire \scs.diff2[7] ;
 wire \scs.diff2[8] ;
 wire \scs.diff2[9] ;
 wire \scs.diff2_d[0] ;
 wire \scs.diff2_d[10] ;
 wire \scs.diff2_d[11] ;
 wire \scs.diff2_d[12] ;
 wire \scs.diff2_d[13] ;
 wire \scs.diff2_d[14] ;
 wire \scs.diff2_d[15] ;
 wire \scs.diff2_d[16] ;
 wire \scs.diff2_d[17] ;
 wire \scs.diff2_d[18] ;
 wire \scs.diff2_d[19] ;
 wire \scs.diff2_d[1] ;
 wire \scs.diff2_d[20] ;
 wire \scs.diff2_d[21] ;
 wire \scs.diff2_d[22] ;
 wire \scs.diff2_d[23] ;
 wire \scs.diff2_d[24] ;
 wire \scs.diff2_d[25] ;
 wire \scs.diff2_d[26] ;
 wire \scs.diff2_d[27] ;
 wire \scs.diff2_d[28] ;
 wire \scs.diff2_d[29] ;
 wire \scs.diff2_d[2] ;
 wire \scs.diff2_d[30] ;
 wire \scs.diff2_d[31] ;
 wire \scs.diff2_d[3] ;
 wire \scs.diff2_d[4] ;
 wire \scs.diff2_d[5] ;
 wire \scs.diff2_d[6] ;
 wire \scs.diff2_d[7] ;
 wire \scs.diff2_d[8] ;
 wire \scs.diff2_d[9] ;
 wire \scs.enable_in ;
 wire \scs.oversample_in[0] ;
 wire \scs.oversample_in[1] ;
 wire \scs.oversample_in[2] ;
 wire \scs.oversample_in[3] ;
 wire \scs.oversample_in[4] ;
 wire \scs.oversample_in[5] ;
 wire \scs.oversample_in[6] ;
 wire \scs.oversample_in[7] ;
 wire \scs.oversample_in[8] ;
 wire \scs.oversample_in[9] ;
 wire \scs.word_count[0] ;
 wire \scs.word_count[1] ;
 wire \scs.word_count[2] ;
 wire \scs.word_count[3] ;
 wire \scs.word_count[4] ;
 wire \scs.word_count[5] ;
 wire \scs.word_count[6] ;
 wire \scs.word_count[7] ;
 wire \scs.word_count[8] ;
 wire \scs.word_count[9] ;
 wire \startup_cnt_reg[0] ;
 wire \startup_cnt_reg[1] ;
 wire \startup_cnt_reg[2] ;

 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__C1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A_N (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A_N (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__C1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__C1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__C1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__C1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__B (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__B (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__A2 (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__C1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__B (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__B (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A_N (.DIODE(_1062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__B (.DIODE(_1062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A1 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__B (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__C1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout572_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout588_A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout591_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout592_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout593_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout600_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold198_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _1729_ (.A(net254),
    .Y(_1447_));
 sky130_fd_sc_hd__inv_2 _1730_ (.A(net428),
    .Y(_1448_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(net255),
    .Y(_1449_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(net258),
    .Y(_1450_));
 sky130_fd_sc_hd__inv_2 _1733_ (.A(net264),
    .Y(_1451_));
 sky130_fd_sc_hd__inv_2 _1734_ (.A(net265),
    .Y(_1452_));
 sky130_fd_sc_hd__inv_2 _1735_ (.A(net267),
    .Y(_1453_));
 sky130_fd_sc_hd__inv_2 _1736_ (.A(net268),
    .Y(_1454_));
 sky130_fd_sc_hd__inv_2 _1737_ (.A(net270),
    .Y(_1455_));
 sky130_fd_sc_hd__inv_2 _1738_ (.A(\scs.diff2_d[27] ),
    .Y(_1456_));
 sky130_fd_sc_hd__inv_2 _1739_ (.A(\scs.diff2[27] ),
    .Y(_1457_));
 sky130_fd_sc_hd__inv_2 _1740_ (.A(net853),
    .Y(_1458_));
 sky130_fd_sc_hd__inv_2 _1741_ (.A(net420),
    .Y(_1459_));
 sky130_fd_sc_hd__inv_2 _1742_ (.A(net833),
    .Y(_1460_));
 sky130_fd_sc_hd__inv_2 _1743_ (.A(net848),
    .Y(_1461_));
 sky130_fd_sc_hd__inv_2 _1744_ (.A(\scs.diff1[27] ),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_2 _1745_ (.A(net659),
    .Y(_1463_));
 sky130_fd_sc_hd__inv_2 _1746_ (.A(net844),
    .Y(_1464_));
 sky130_fd_sc_hd__inv_2 _1747_ (.A(net414),
    .Y(_1465_));
 sky130_fd_sc_hd__inv_2 _1748_ (.A(net825),
    .Y(_1466_));
 sky130_fd_sc_hd__inv_2 _1749_ (.A(net823),
    .Y(_1467_));
 sky130_fd_sc_hd__inv_2 _1750_ (.A(net775),
    .Y(_1468_));
 sky130_fd_sc_hd__inv_2 _1751_ (.A(net809),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _1752_ (.A(net651),
    .Y(_1470_));
 sky130_fd_sc_hd__inv_2 _1753_ (.A(net308),
    .Y(_1471_));
 sky130_fd_sc_hd__inv_2 _1754_ (.A(net311),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _1755_ (.A(net325),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _1756_ (.A(net333),
    .Y(_1474_));
 sky130_fd_sc_hd__inv_2 _1757_ (.A(\scs.acc2[31] ),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _1758_ (.A(\scs.acc3_d2[6] ),
    .Y(_1476_));
 sky130_fd_sc_hd__inv_2 _1759_ (.A(net706),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_2 _1760_ (.A(net581),
    .Y(_1478_));
 sky130_fd_sc_hd__inv_2 _1761_ (.A(\scs.oversample_in[1] ),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _1762_ (.A(\scs.oversample_in[2] ),
    .Y(_1480_));
 sky130_fd_sc_hd__inv_2 _1763_ (.A(\scs.oversample_in[3] ),
    .Y(_1481_));
 sky130_fd_sc_hd__inv_2 _1764_ (.A(\scs.oversample_in[6] ),
    .Y(_1482_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(\scs.oversample_in[8] ),
    .Y(_1483_));
 sky130_fd_sc_hd__inv_2 _1766_ (.A(\scs.oversample_in[9] ),
    .Y(_1484_));
 sky130_fd_sc_hd__inv_2 _1767_ (.A(\scs.oversample_in[0] ),
    .Y(_1485_));
 sky130_fd_sc_hd__and2_1 _1768_ (.A(\scs.data_valid_out ),
    .B(output_en_reg),
    .X(net56));
 sky130_fd_sc_hd__or3b_1 _1769_ (.A(net472),
    .B(net805),
    .C_N(net840),
    .X(_1486_));
 sky130_fd_sc_hd__nand3_1 _1770_ (.A(net425),
    .B(\scs.data_valid_out ),
    .C(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(net425),
    .B(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(_1487_),
    .A1(_1488_),
    .S(net863),
    .X(_1489_));
 sky130_fd_sc_hd__nor2_1 _1773_ (.A(net575),
    .B(_1489_),
    .Y(_0000_));
 sky130_fd_sc_hd__a31o_1 _1774_ (.A1(net472),
    .A2(net805),
    .A3(\scs.data_valid_out ),
    .B1(net236),
    .X(_1490_));
 sky130_fd_sc_hd__inv_2 _1775_ (.A(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__and4b_1 _1776_ (.A_N(\startup_cnt_reg[1] ),
    .B(net805),
    .C(\scs.data_valid_out ),
    .D(net426),
    .X(_1492_));
 sky130_fd_sc_hd__a21oi_1 _1777_ (.A1(net472),
    .A2(_1491_),
    .B1(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__nor2_1 _1778_ (.A(net575),
    .B(_1493_),
    .Y(_0001_));
 sky130_fd_sc_hd__nand3b_1 _1779_ (.A_N(net857),
    .B(net472),
    .C(net805),
    .Y(_1494_));
 sky130_fd_sc_hd__o2bb2a_1 _1780_ (.A1_N(net840),
    .A2_N(_1491_),
    .B1(_1494_),
    .B2(_1487_),
    .X(_1495_));
 sky130_fd_sc_hd__nor2_1 _1781_ (.A(net576),
    .B(_1495_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_1 _1782_ (.A(net636),
    .B(net509),
    .X(_0003_));
 sky130_fd_sc_hd__nor3_1 _1783_ (.A(net236),
    .B(net575),
    .C(net841),
    .Y(_0004_));
 sky130_fd_sc_hd__or2_1 _1784_ (.A(net574),
    .B(net2),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _1785_ (.A(net575),
    .B(net3),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _1786_ (.A(net576),
    .B(net4),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _1787_ (.A(net581),
    .B(net5),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _1788_ (.A(net580),
    .B(net6),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _1789_ (.A(net580),
    .B(net7),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _1790_ (.A(net580),
    .B(net8),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1791_ (.A(net580),
    .B(net9),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _1792_ (.A(net511),
    .B(net10),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _1793_ (.A(net511),
    .B(net11),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1794_ (.A(net483),
    .B(net1),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _1795_ (.A(net425),
    .B(\scs.decimation_en ),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _1796_ (.A(net425),
    .B(\scs.decimation_en ),
    .Y(_1497_));
 sky130_fd_sc_hd__and2b_1 _1797_ (.A_N(\scs.diff1_d[0] ),
    .B(\scs.diff1[0] ),
    .X(_1498_));
 sky130_fd_sc_hd__nand2b_1 _1798_ (.A_N(\scs.diff1[0] ),
    .B(\scs.diff1_d[0] ),
    .Y(_1499_));
 sky130_fd_sc_hd__or3b_1 _1799_ (.A(net74),
    .B(_1498_),
    .C_N(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__o211a_1 _1800_ (.A1(net750),
    .A2(net153),
    .B1(_1500_),
    .C1(net475),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _1801_ (.A_N(\scs.diff1_d[1] ),
    .B(\scs.diff1[1] ),
    .X(_1501_));
 sky130_fd_sc_hd__nand2b_1 _1802_ (.A_N(\scs.diff1[1] ),
    .B(\scs.diff1_d[1] ),
    .Y(_1502_));
 sky130_fd_sc_hd__and2b_1 _1803_ (.A_N(_1501_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__xnor2_1 _1804_ (.A(_1499_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(net153),
    .B(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__o211a_1 _1806_ (.A1(net699),
    .A2(net153),
    .B1(_1505_),
    .C1(net476),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_2 _1807_ (.A1(_1499_),
    .A2(_1502_),
    .B1(_1501_),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2b_1 _1808_ (.A_N(\scs.diff1[2] ),
    .B(\scs.diff1_d[2] ),
    .Y(_1507_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2b_1 _1810_ (.A_N(\scs.diff1_d[2] ),
    .B(\scs.diff1[2] ),
    .Y(_1509_));
 sky130_fd_sc_hd__a21oi_1 _1811_ (.A1(_1507_),
    .A2(_1509_),
    .B1(_1506_),
    .Y(_1510_));
 sky130_fd_sc_hd__a31o_1 _1812_ (.A1(_1506_),
    .A2(_1507_),
    .A3(_1509_),
    .B1(net73),
    .X(_1511_));
 sky130_fd_sc_hd__o221a_1 _1813_ (.A1(net735),
    .A2(net154),
    .B1(_1510_),
    .B2(_1511_),
    .C1(net475),
    .X(_0018_));
 sky130_fd_sc_hd__o21ai_2 _1814_ (.A1(_1506_),
    .A2(_1508_),
    .B1(_1509_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2b_1 _1815_ (.A_N(\scs.diff1[3] ),
    .B(\scs.diff1_d[3] ),
    .Y(_1513_));
 sky130_fd_sc_hd__inv_2 _1816_ (.A(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__and2b_1 _1817_ (.A_N(\scs.diff1_d[3] ),
    .B(\scs.diff1[3] ),
    .X(_1515_));
 sky130_fd_sc_hd__o21a_1 _1818_ (.A1(_1514_),
    .A2(_1515_),
    .B1(_1512_),
    .X(_1516_));
 sky130_fd_sc_hd__o31ai_1 _1819_ (.A1(_1512_),
    .A2(_1514_),
    .A3(_1515_),
    .B1(net155),
    .Y(_1517_));
 sky130_fd_sc_hd__o221a_1 _1820_ (.A1(net756),
    .A2(net154),
    .B1(_1516_),
    .B2(_1517_),
    .C1(net475),
    .X(_0019_));
 sky130_fd_sc_hd__a21o_1 _1821_ (.A1(_1512_),
    .A2(_1513_),
    .B1(_1515_),
    .X(_1518_));
 sky130_fd_sc_hd__and2b_1 _1822_ (.A_N(\scs.diff1_d[4] ),
    .B(\scs.diff1[4] ),
    .X(_1519_));
 sky130_fd_sc_hd__and2b_1 _1823_ (.A_N(\scs.diff1[4] ),
    .B(\scs.diff1_d[4] ),
    .X(_1520_));
 sky130_fd_sc_hd__nor2_1 _1824_ (.A(_1519_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__xor2_1 _1825_ (.A(_1518_),
    .B(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__or2_1 _1826_ (.A(net672),
    .B(net158),
    .X(_1523_));
 sky130_fd_sc_hd__o211a_1 _1827_ (.A1(net77),
    .A2(_1522_),
    .B1(_1523_),
    .C1(net480),
    .X(_0020_));
 sky130_fd_sc_hd__nand2b_1 _1828_ (.A_N(\scs.diff1[5] ),
    .B(\scs.diff1_d[5] ),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2b_1 _1829_ (.A_N(\scs.diff1_d[5] ),
    .B(\scs.diff1[5] ),
    .Y(_1525_));
 sky130_fd_sc_hd__nand2_1 _1830_ (.A(_1524_),
    .B(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__inv_2 _1831_ (.A(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__a21o_1 _1832_ (.A1(_1518_),
    .A2(_1521_),
    .B1(_1519_),
    .X(_1528_));
 sky130_fd_sc_hd__nor2_1 _1833_ (.A(_1526_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a21o_1 _1834_ (.A1(_1526_),
    .A2(_1528_),
    .B1(net77),
    .X(_1530_));
 sky130_fd_sc_hd__o221a_1 _1835_ (.A1(net722),
    .A2(net158),
    .B1(_1529_),
    .B2(_1530_),
    .C1(net480),
    .X(_0021_));
 sky130_fd_sc_hd__a21bo_1 _1836_ (.A1(_1519_),
    .A2(_1524_),
    .B1_N(_1525_),
    .X(_1531_));
 sky130_fd_sc_hd__a31o_1 _1837_ (.A1(_1518_),
    .A2(_1521_),
    .A3(_1527_),
    .B1(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__and2b_1 _1838_ (.A_N(\scs.diff1_d[6] ),
    .B(\scs.diff1[6] ),
    .X(_1533_));
 sky130_fd_sc_hd__and2b_1 _1839_ (.A_N(\scs.diff1[6] ),
    .B(\scs.diff1_d[6] ),
    .X(_1534_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(_1533_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__nand2_1 _1841_ (.A(_1532_),
    .B(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__or2_1 _1842_ (.A(_1532_),
    .B(_1535_),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_1 _1843_ (.A1(_1536_),
    .A2(_1537_),
    .B1(net77),
    .X(_1538_));
 sky130_fd_sc_hd__o211a_1 _1844_ (.A1(net697),
    .A2(net159),
    .B1(_1538_),
    .C1(net481),
    .X(_0022_));
 sky130_fd_sc_hd__nand2b_1 _1845_ (.A_N(net418),
    .B(\scs.diff1_d[7] ),
    .Y(_1539_));
 sky130_fd_sc_hd__and2b_1 _1846_ (.A_N(\scs.diff1_d[7] ),
    .B(net418),
    .X(_1540_));
 sky130_fd_sc_hd__nand2b_1 _1847_ (.A_N(\scs.diff1_d[7] ),
    .B(net418),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _1848_ (.A(_1539_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__a21o_1 _1849_ (.A1(_1532_),
    .A2(_1535_),
    .B1(_1533_),
    .X(_1543_));
 sky130_fd_sc_hd__nor2_1 _1850_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__a21o_1 _1851_ (.A1(_1542_),
    .A2(_1543_),
    .B1(net78),
    .X(_1545_));
 sky130_fd_sc_hd__o221a_1 _1852_ (.A1(net657),
    .A2(net158),
    .B1(_1544_),
    .B2(_1545_),
    .C1(net481),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _1853_ (.A(_1533_),
    .B(_1539_),
    .X(_1546_));
 sky130_fd_sc_hd__a311o_1 _1854_ (.A1(_1532_),
    .A2(_1535_),
    .A3(_1539_),
    .B1(_1540_),
    .C1(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__and2b_1 _1855_ (.A_N(\scs.diff1_d[8] ),
    .B(\scs.diff1[8] ),
    .X(_1548_));
 sky130_fd_sc_hd__and2b_1 _1856_ (.A_N(\scs.diff1[8] ),
    .B(\scs.diff1_d[8] ),
    .X(_1549_));
 sky130_fd_sc_hd__nor2_1 _1857_ (.A(_1548_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__xor2_1 _1858_ (.A(_1547_),
    .B(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__or2_1 _1859_ (.A(net680),
    .B(net173),
    .X(_1552_));
 sky130_fd_sc_hd__o211a_1 _1860_ (.A1(net90),
    .A2(_1551_),
    .B1(_1552_),
    .C1(net494),
    .X(_0024_));
 sky130_fd_sc_hd__nand2b_1 _1861_ (.A_N(\scs.diff1[9] ),
    .B(\scs.diff1_d[9] ),
    .Y(_1553_));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__and2b_1 _1863_ (.A_N(\scs.diff1_d[9] ),
    .B(\scs.diff1[9] ),
    .X(_1555_));
 sky130_fd_sc_hd__nor2_1 _1864_ (.A(_1554_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__a21oi_1 _1865_ (.A1(_1547_),
    .A2(_1550_),
    .B1(_1548_),
    .Y(_1557_));
 sky130_fd_sc_hd__and2_1 _1866_ (.A(_1556_),
    .B(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__o21ai_1 _1867_ (.A1(_1556_),
    .A2(_1557_),
    .B1(net173),
    .Y(_1559_));
 sky130_fd_sc_hd__o221a_1 _1868_ (.A1(net728),
    .A2(net173),
    .B1(_1558_),
    .B2(_1559_),
    .C1(net493),
    .X(_0025_));
 sky130_fd_sc_hd__nand2b_1 _1869_ (.A_N(\scs.diff1_d[10] ),
    .B(\scs.diff1[10] ),
    .Y(_1560_));
 sky130_fd_sc_hd__inv_2 _1870_ (.A(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2b_1 _1871_ (.A_N(\scs.diff1[10] ),
    .B(\scs.diff1_d[10] ),
    .Y(_1562_));
 sky130_fd_sc_hd__a211o_1 _1872_ (.A1(_1547_),
    .A2(_1550_),
    .B1(_1555_),
    .C1(_1548_),
    .X(_1563_));
 sky130_fd_sc_hd__a22oi_1 _1873_ (.A1(_1560_),
    .A2(_1562_),
    .B1(_1563_),
    .B2(_1553_),
    .Y(_1564_));
 sky130_fd_sc_hd__a41o_1 _1874_ (.A1(_1553_),
    .A2(_1560_),
    .A3(_1562_),
    .A4(_1563_),
    .B1(net90),
    .X(_1565_));
 sky130_fd_sc_hd__o2bb2a_1 _1875_ (.A1_N(net691),
    .A2_N(net91),
    .B1(_1564_),
    .B2(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(net574),
    .B(_1566_),
    .Y(_0026_));
 sky130_fd_sc_hd__and2b_1 _1877_ (.A_N(\scs.diff1_d[11] ),
    .B(\scs.diff1[11] ),
    .X(_1567_));
 sky130_fd_sc_hd__nand2b_1 _1878_ (.A_N(\scs.diff1[11] ),
    .B(\scs.diff1_d[11] ),
    .Y(_1568_));
 sky130_fd_sc_hd__nand2b_1 _1879_ (.A_N(_1567_),
    .B(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__a31o_1 _1880_ (.A1(_1553_),
    .A2(_1562_),
    .A3(_1563_),
    .B1(_1561_),
    .X(_1570_));
 sky130_fd_sc_hd__xnor2_1 _1881_ (.A(_1569_),
    .B(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(net674),
    .A1(_1571_),
    .S(net174),
    .X(_1572_));
 sky130_fd_sc_hd__and2_1 _1883_ (.A(net493),
    .B(_1572_),
    .X(_0027_));
 sky130_fd_sc_hd__a21oi_2 _1884_ (.A1(_1568_),
    .A2(_1570_),
    .B1(_1567_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2b_1 _1885_ (.A_N(\scs.diff1_d[12] ),
    .B(\scs.diff1[12] ),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2b_1 _1886_ (.A_N(\scs.diff1[12] ),
    .B(\scs.diff1_d[12] ),
    .Y(_1575_));
 sky130_fd_sc_hd__nand2_1 _1887_ (.A(_1574_),
    .B(_1575_),
    .Y(_1576_));
 sky130_fd_sc_hd__or2_1 _1888_ (.A(_1573_),
    .B(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__xnor2_1 _1889_ (.A(_1573_),
    .B(_1576_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _1890_ (.A(net178),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__o211a_1 _1891_ (.A1(net733),
    .A2(net178),
    .B1(_1579_),
    .C1(net498),
    .X(_0028_));
 sky130_fd_sc_hd__and2b_1 _1892_ (.A_N(\scs.diff1[13] ),
    .B(\scs.diff1_d[13] ),
    .X(_1580_));
 sky130_fd_sc_hd__nand2b_1 _1893_ (.A_N(\scs.diff1_d[13] ),
    .B(\scs.diff1[13] ),
    .Y(_1581_));
 sky130_fd_sc_hd__and2b_1 _1894_ (.A_N(_1580_),
    .B(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__inv_2 _1895_ (.A(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__a21oi_1 _1896_ (.A1(_1574_),
    .A2(_1577_),
    .B1(_1582_),
    .Y(_1584_));
 sky130_fd_sc_hd__a31o_1 _1897_ (.A1(_1574_),
    .A2(_1577_),
    .A3(_1582_),
    .B1(net94),
    .X(_1585_));
 sky130_fd_sc_hd__o221a_1 _1898_ (.A1(net763),
    .A2(net178),
    .B1(_1584_),
    .B2(_1585_),
    .C1(net498),
    .X(_0029_));
 sky130_fd_sc_hd__nand2b_1 _1899_ (.A_N(\scs.diff1_d[14] ),
    .B(\scs.diff1[14] ),
    .Y(_1586_));
 sky130_fd_sc_hd__nand2b_1 _1900_ (.A_N(\scs.diff1[14] ),
    .B(\scs.diff1_d[14] ),
    .Y(_1587_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_1586_),
    .B(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__or2_1 _1902_ (.A(_1574_),
    .B(_1580_),
    .X(_1589_));
 sky130_fd_sc_hd__o311a_1 _1903_ (.A1(_1573_),
    .A2(_1576_),
    .A3(_1583_),
    .B1(_1589_),
    .C1(_1581_),
    .X(_1590_));
 sky130_fd_sc_hd__or2_1 _1904_ (.A(_1588_),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__xor2_1 _1905_ (.A(_1588_),
    .B(_1590_),
    .X(_1592_));
 sky130_fd_sc_hd__or2_1 _1906_ (.A(net621),
    .B(net179),
    .X(_1593_));
 sky130_fd_sc_hd__o211a_1 _1907_ (.A1(net94),
    .A2(_1592_),
    .B1(_1593_),
    .C1(net524),
    .X(_0030_));
 sky130_fd_sc_hd__xnor2_2 _1908_ (.A(\scs.diff1_d[15] ),
    .B(net417),
    .Y(_1594_));
 sky130_fd_sc_hd__inv_2 _1909_ (.A(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__a21oi_1 _1910_ (.A1(_1586_),
    .A2(_1591_),
    .B1(_1594_),
    .Y(_1596_));
 sky130_fd_sc_hd__a31o_1 _1911_ (.A1(_1586_),
    .A2(_1591_),
    .A3(_1594_),
    .B1(net95),
    .X(_1597_));
 sky130_fd_sc_hd__o221a_1 _1912_ (.A1(net667),
    .A2(net179),
    .B1(_1596_),
    .B2(_1597_),
    .C1(net497),
    .X(_0031_));
 sky130_fd_sc_hd__nand2b_1 _1913_ (.A_N(\scs.diff1_d[16] ),
    .B(\scs.diff1[16] ),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2b_1 _1914_ (.A_N(\scs.diff1[16] ),
    .B(\scs.diff1_d[16] ),
    .Y(_1599_));
 sky130_fd_sc_hd__nand2_1 _1915_ (.A(_1598_),
    .B(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__o21ba_1 _1916_ (.A1(_1466_),
    .A2(net417),
    .B1_N(_1586_),
    .X(_1601_));
 sky130_fd_sc_hd__a21oi_1 _1917_ (.A1(_1466_),
    .A2(net417),
    .B1(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__o31a_1 _1918_ (.A1(_1588_),
    .A2(_1590_),
    .A3(_1595_),
    .B1(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__or2_1 _1919_ (.A(_1600_),
    .B(net66),
    .X(_1604_));
 sky130_fd_sc_hd__nand2_1 _1920_ (.A(_1600_),
    .B(net66),
    .Y(_1605_));
 sky130_fd_sc_hd__a21o_1 _1921_ (.A1(_1604_),
    .A2(_1605_),
    .B1(net110),
    .X(_1606_));
 sky130_fd_sc_hd__o211a_1 _1922_ (.A1(net724),
    .A2(net195),
    .B1(_1606_),
    .C1(net525),
    .X(_0032_));
 sky130_fd_sc_hd__and2b_1 _1923_ (.A_N(\scs.diff1_d[17] ),
    .B(net416),
    .X(_1607_));
 sky130_fd_sc_hd__nand2b_1 _1924_ (.A_N(\scs.diff1_d[17] ),
    .B(net416),
    .Y(_1608_));
 sky130_fd_sc_hd__and2b_1 _1925_ (.A_N(net416),
    .B(\scs.diff1_d[17] ),
    .X(_1609_));
 sky130_fd_sc_hd__nor2_1 _1926_ (.A(_1607_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21a_1 _1927_ (.A1(_1600_),
    .A2(net66),
    .B1(_1598_),
    .X(_1611_));
 sky130_fd_sc_hd__xnor2_1 _1928_ (.A(_1610_),
    .B(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__or2_1 _1929_ (.A(net770),
    .B(net195),
    .X(_1613_));
 sky130_fd_sc_hd__o211a_1 _1930_ (.A1(net110),
    .A2(_1612_),
    .B1(_1613_),
    .C1(net524),
    .X(_0033_));
 sky130_fd_sc_hd__nand2b_1 _1931_ (.A_N(\scs.diff1_d[18] ),
    .B(net415),
    .Y(_1614_));
 sky130_fd_sc_hd__xnor2_2 _1932_ (.A(\scs.diff1_d[18] ),
    .B(net415),
    .Y(_1615_));
 sky130_fd_sc_hd__inv_2 _1933_ (.A(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__a21o_1 _1934_ (.A1(_1608_),
    .A2(_1611_),
    .B1(_1609_),
    .X(_1617_));
 sky130_fd_sc_hd__or2_1 _1935_ (.A(_1616_),
    .B(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__xnor2_1 _1936_ (.A(_1615_),
    .B(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__or2_1 _1937_ (.A(net762),
    .B(net196),
    .X(_1620_));
 sky130_fd_sc_hd__o211a_1 _1938_ (.A1(net110),
    .A2(_1619_),
    .B1(_1620_),
    .C1(net527),
    .X(_0034_));
 sky130_fd_sc_hd__xnor2_1 _1939_ (.A(\scs.diff1_d[19] ),
    .B(net414),
    .Y(_1621_));
 sky130_fd_sc_hd__a21oi_1 _1940_ (.A1(_1614_),
    .A2(_1618_),
    .B1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__a31o_1 _1941_ (.A1(_1614_),
    .A2(_1618_),
    .A3(_1621_),
    .B1(net111),
    .X(_1623_));
 sky130_fd_sc_hd__o221a_1 _1942_ (.A1(net639),
    .A2(net195),
    .B1(_1622_),
    .B2(_1623_),
    .C1(net524),
    .X(_0035_));
 sky130_fd_sc_hd__and2b_1 _1943_ (.A_N(\scs.diff1_d[20] ),
    .B(\scs.diff1[20] ),
    .X(_1624_));
 sky130_fd_sc_hd__and2b_1 _1944_ (.A_N(\scs.diff1[20] ),
    .B(\scs.diff1_d[20] ),
    .X(_1625_));
 sky130_fd_sc_hd__nor2_1 _1945_ (.A(_1624_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__nand2_1 _1946_ (.A(_1615_),
    .B(_1621_),
    .Y(_1627_));
 sky130_fd_sc_hd__a211o_1 _1947_ (.A1(_1598_),
    .A2(_1608_),
    .B1(_1609_),
    .C1(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__o21ai_1 _1948_ (.A1(_1464_),
    .A2(net414),
    .B1(net415),
    .Y(_1629_));
 sky130_fd_sc_hd__o221a_1 _1949_ (.A1(\scs.diff1_d[19] ),
    .A2(_1465_),
    .B1(\scs.diff1_d[18] ),
    .B2(_1629_),
    .C1(_1628_),
    .X(_1630_));
 sky130_fd_sc_hd__or4_1 _1950_ (.A(_1600_),
    .B(_1607_),
    .C(_1609_),
    .D(_1627_),
    .X(_1631_));
 sky130_fd_sc_hd__o21ai_1 _1951_ (.A1(net66),
    .A2(_1631_),
    .B1(_1630_),
    .Y(_1632_));
 sky130_fd_sc_hd__xnor2_1 _1952_ (.A(_1626_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__nor2_1 _1953_ (.A(net718),
    .B(net199),
    .Y(_1634_));
 sky130_fd_sc_hd__a211oi_1 _1954_ (.A1(net199),
    .A2(_1633_),
    .B1(_1634_),
    .C1(net593),
    .Y(_0036_));
 sky130_fd_sc_hd__and2b_1 _1955_ (.A_N(\scs.diff1_d[21] ),
    .B(net413),
    .X(_1635_));
 sky130_fd_sc_hd__nand2b_1 _1956_ (.A_N(\scs.diff1_d[21] ),
    .B(net413),
    .Y(_1636_));
 sky130_fd_sc_hd__and2b_1 _1957_ (.A_N(net413),
    .B(\scs.diff1_d[21] ),
    .X(_1637_));
 sky130_fd_sc_hd__nor2_1 _1958_ (.A(_1635_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a21oi_1 _1959_ (.A1(_1626_),
    .A2(_1632_),
    .B1(_1624_),
    .Y(_1639_));
 sky130_fd_sc_hd__and2_1 _1960_ (.A(_1638_),
    .B(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__o21ai_1 _1961_ (.A1(_1638_),
    .A2(_1639_),
    .B1(net199),
    .Y(_1641_));
 sky130_fd_sc_hd__o221a_1 _1962_ (.A1(net650),
    .A2(net200),
    .B1(_1640_),
    .B2(_1641_),
    .C1(net527),
    .X(_0037_));
 sky130_fd_sc_hd__nand2b_1 _1963_ (.A_N(\scs.diff1_d[22] ),
    .B(\scs.diff1[22] ),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2b_1 _1964_ (.A_N(\scs.diff1[22] ),
    .B(\scs.diff1_d[22] ),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(_1642_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__a21o_1 _1966_ (.A1(_1636_),
    .A2(_1639_),
    .B1(_1637_),
    .X(_1645_));
 sky130_fd_sc_hd__nand2_1 _1967_ (.A(_1644_),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__or2_1 _1968_ (.A(_1644_),
    .B(_1645_),
    .X(_1647_));
 sky130_fd_sc_hd__a21o_1 _1969_ (.A1(_1646_),
    .A2(_1647_),
    .B1(net113),
    .X(_1648_));
 sky130_fd_sc_hd__o211a_1 _1970_ (.A1(net785),
    .A2(net200),
    .B1(_1648_),
    .C1(net538),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _1971_ (.A(\scs.diff1_d[23] ),
    .B(_1463_),
    .X(_1649_));
 sky130_fd_sc_hd__or2_1 _1972_ (.A(\scs.diff1_d[23] ),
    .B(_1463_),
    .X(_1650_));
 sky130_fd_sc_hd__and2b_1 _1973_ (.A_N(_1649_),
    .B(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__a21oi_1 _1974_ (.A1(_1642_),
    .A2(_1647_),
    .B1(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__and3_1 _1975_ (.A(_1642_),
    .B(_1647_),
    .C(_1651_),
    .X(_1653_));
 sky130_fd_sc_hd__or2_1 _1976_ (.A(net684),
    .B(net216),
    .X(_1654_));
 sky130_fd_sc_hd__o311a_1 _1977_ (.A1(net126),
    .A2(_1652_),
    .A3(_1653_),
    .B1(_1654_),
    .C1(net538),
    .X(_0039_));
 sky130_fd_sc_hd__nand2b_1 _1978_ (.A_N(\scs.diff1_d[24] ),
    .B(\scs.diff1[24] ),
    .Y(_1655_));
 sky130_fd_sc_hd__nand2b_1 _1979_ (.A_N(\scs.diff1[24] ),
    .B(\scs.diff1_d[24] ),
    .Y(_1656_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(_1655_),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2b_1 _1981_ (.A_N(_1644_),
    .B(_1651_),
    .Y(_1658_));
 sky130_fd_sc_hd__or4b_1 _1982_ (.A(_1635_),
    .B(_1637_),
    .C(_1658_),
    .D_N(_1626_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2b_1 _1983_ (.A_N(_1637_),
    .B(_1624_),
    .Y(_1660_));
 sky130_fd_sc_hd__a21o_1 _1984_ (.A1(_1636_),
    .A2(_1660_),
    .B1(_1658_),
    .X(_1661_));
 sky130_fd_sc_hd__a21o_1 _1985_ (.A1(_1642_),
    .A2(_1650_),
    .B1(_1649_),
    .X(_1662_));
 sky130_fd_sc_hd__o211a_1 _1986_ (.A1(_1630_),
    .A2(_1659_),
    .B1(_1661_),
    .C1(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__o31a_1 _1987_ (.A1(_1603_),
    .A2(_1631_),
    .A3(_1659_),
    .B1(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__or2_1 _1988_ (.A(_1657_),
    .B(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__nand2_1 _1989_ (.A(_1657_),
    .B(_1664_),
    .Y(_1666_));
 sky130_fd_sc_hd__a21o_1 _1990_ (.A1(_1665_),
    .A2(_1666_),
    .B1(net126),
    .X(_1667_));
 sky130_fd_sc_hd__o211a_1 _1991_ (.A1(net740),
    .A2(net216),
    .B1(_1667_),
    .C1(net538),
    .X(_0040_));
 sky130_fd_sc_hd__nand2b_1 _1992_ (.A_N(\scs.diff1_d[25] ),
    .B(\scs.diff1[25] ),
    .Y(_1668_));
 sky130_fd_sc_hd__and2b_1 _1993_ (.A_N(\scs.diff1[25] ),
    .B(\scs.diff1_d[25] ),
    .X(_1669_));
 sky130_fd_sc_hd__inv_2 _1994_ (.A(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(_1668_),
    .B(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__nand2_1 _1996_ (.A(_1655_),
    .B(_1665_),
    .Y(_1672_));
 sky130_fd_sc_hd__xnor2_1 _1997_ (.A(_1671_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__or2_1 _1998_ (.A(net713),
    .B(net215),
    .X(_1674_));
 sky130_fd_sc_hd__o211a_1 _1999_ (.A1(net125),
    .A2(_1673_),
    .B1(_1674_),
    .C1(net539),
    .X(_0041_));
 sky130_fd_sc_hd__nand2b_1 _2000_ (.A_N(\scs.diff1_d[26] ),
    .B(\scs.diff1[26] ),
    .Y(_1675_));
 sky130_fd_sc_hd__xnor2_2 _2001_ (.A(\scs.diff1_d[26] ),
    .B(\scs.diff1[26] ),
    .Y(_1676_));
 sky130_fd_sc_hd__inv_2 _2002_ (.A(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__a31o_1 _2003_ (.A1(_1655_),
    .A2(_1665_),
    .A3(_1668_),
    .B1(_1669_),
    .X(_1678_));
 sky130_fd_sc_hd__or2_1 _2004_ (.A(_1677_),
    .B(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__xnor2_1 _2005_ (.A(_1676_),
    .B(_1678_),
    .Y(_1680_));
 sky130_fd_sc_hd__or2_1 _2006_ (.A(\scs.diff2[26] ),
    .B(net215),
    .X(_1681_));
 sky130_fd_sc_hd__o211a_1 _2007_ (.A1(net125),
    .A2(_1680_),
    .B1(_1681_),
    .C1(net543),
    .X(_0042_));
 sky130_fd_sc_hd__xnor2_1 _2008_ (.A(\scs.diff1_d[27] ),
    .B(\scs.diff1[27] ),
    .Y(_1682_));
 sky130_fd_sc_hd__a21oi_1 _2009_ (.A1(_1675_),
    .A2(_1679_),
    .B1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__a31o_1 _2010_ (.A1(_1675_),
    .A2(_1679_),
    .A3(_1682_),
    .B1(net131),
    .X(_1684_));
 sky130_fd_sc_hd__o221a_1 _2011_ (.A1(net846),
    .A2(net219),
    .B1(_1683_),
    .B2(_1684_),
    .C1(net543),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_1 _2012_ (.A(_1676_),
    .B(_1682_),
    .Y(_1685_));
 sky130_fd_sc_hd__or4_1 _2013_ (.A(_1657_),
    .B(_1664_),
    .C(_1671_),
    .D(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__a211o_1 _2014_ (.A1(_1655_),
    .A2(_1668_),
    .B1(_1669_),
    .C1(_1685_),
    .X(_1687_));
 sky130_fd_sc_hd__a21o_1 _2015_ (.A1(\scs.diff1_d[27] ),
    .A2(_1462_),
    .B1(_1675_),
    .X(_1688_));
 sky130_fd_sc_hd__o2111a_1 _2016_ (.A1(\scs.diff1_d[27] ),
    .A2(_1462_),
    .B1(_1686_),
    .C1(_1687_),
    .D1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__and2b_1 _2017_ (.A_N(\scs.diff1[28] ),
    .B(\scs.diff1_d[28] ),
    .X(_1690_));
 sky130_fd_sc_hd__nand2b_1 _2018_ (.A_N(\scs.diff1_d[28] ),
    .B(\scs.diff1[28] ),
    .Y(_1691_));
 sky130_fd_sc_hd__and2b_1 _2019_ (.A_N(_1690_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__and2_1 _2020_ (.A(_1689_),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__o21ai_1 _2021_ (.A1(_1689_),
    .A2(_1692_),
    .B1(net219),
    .Y(_1694_));
 sky130_fd_sc_hd__o221a_1 _2022_ (.A1(net744),
    .A2(net219),
    .B1(_1693_),
    .B2(_1694_),
    .C1(net543),
    .X(_0044_));
 sky130_fd_sc_hd__o21ai_2 _2023_ (.A1(_1689_),
    .A2(_1690_),
    .B1(_1691_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2b_1 _2024_ (.A_N(\scs.diff1[29] ),
    .B(\scs.diff1_d[29] ),
    .Y(_1696_));
 sky130_fd_sc_hd__and2b_1 _2025_ (.A_N(\scs.diff1_d[29] ),
    .B(\scs.diff1[29] ),
    .X(_1697_));
 sky130_fd_sc_hd__inv_2 _2026_ (.A(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _2027_ (.A(_1696_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _2028_ (.A(_1695_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__a21o_1 _2029_ (.A1(_1695_),
    .A2(_1699_),
    .B1(net132),
    .X(_1701_));
 sky130_fd_sc_hd__o221a_1 _2030_ (.A1(net783),
    .A2(net220),
    .B1(_1700_),
    .B2(_1701_),
    .C1(net544),
    .X(_0045_));
 sky130_fd_sc_hd__nand2b_1 _2031_ (.A_N(\scs.diff1_d[30] ),
    .B(\scs.diff1[30] ),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2b_1 _2032_ (.A_N(\scs.diff1[30] ),
    .B(\scs.diff1_d[30] ),
    .Y(_1703_));
 sky130_fd_sc_hd__a21o_1 _2033_ (.A1(_1695_),
    .A2(_1696_),
    .B1(_1697_),
    .X(_1704_));
 sky130_fd_sc_hd__a21o_1 _2034_ (.A1(_1702_),
    .A2(_1703_),
    .B1(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__a31oi_1 _2035_ (.A1(_1702_),
    .A2(_1703_),
    .A3(_1704_),
    .B1(net138),
    .Y(_1706_));
 sky130_fd_sc_hd__a22o_1 _2036_ (.A1(net777),
    .A2(net138),
    .B1(_1705_),
    .B2(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__and2_1 _2037_ (.A(net550),
    .B(_1707_),
    .X(_0046_));
 sky130_fd_sc_hd__a21bo_1 _2038_ (.A1(_1703_),
    .A2(_1704_),
    .B1_N(_1702_),
    .X(_1708_));
 sky130_fd_sc_hd__xor2_1 _2039_ (.A(\scs.diff1_d[31] ),
    .B(\scs.diff1[31] ),
    .X(_1709_));
 sky130_fd_sc_hd__xnor2_1 _2040_ (.A(_1708_),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__or2_1 _2041_ (.A(net707),
    .B(net220),
    .X(_1711_));
 sky130_fd_sc_hd__o211a_1 _2042_ (.A1(net131),
    .A2(_1710_),
    .B1(_1711_),
    .C1(net544),
    .X(_0047_));
 sky130_fd_sc_hd__nand2b_1 _2043_ (.A_N(net361),
    .B(\scs.acc3_d2[0] ),
    .Y(_1712_));
 sky130_fd_sc_hd__and2b_1 _2044_ (.A_N(net789),
    .B(net361),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_1 _2045_ (.A(net163),
    .B(net696),
    .Y(_1714_));
 sky130_fd_sc_hd__o221a_1 _2046_ (.A1(net751),
    .A2(net163),
    .B1(_1713_),
    .B2(_1714_),
    .C1(net489),
    .X(_0048_));
 sky130_fd_sc_hd__and2b_1 _2047_ (.A_N(\scs.acc3_d2[1] ),
    .B(net359),
    .X(_1715_));
 sky130_fd_sc_hd__nand2b_1 _2048_ (.A_N(net359),
    .B(\scs.acc3_d2[1] ),
    .Y(_1716_));
 sky130_fd_sc_hd__and2b_1 _2049_ (.A_N(_1715_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__xnor2_1 _2050_ (.A(_1712_),
    .B(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__nand2_1 _2051_ (.A(net161),
    .B(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__o211a_1 _2052_ (.A1(net693),
    .A2(net161),
    .B1(_1719_),
    .C1(net484),
    .X(_0049_));
 sky130_fd_sc_hd__a21oi_1 _2053_ (.A1(_1712_),
    .A2(_1716_),
    .B1(_1715_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2b_1 _2054_ (.A_N(net358),
    .B(\scs.acc3_d2[2] ),
    .Y(_1721_));
 sky130_fd_sc_hd__inv_2 _2055_ (.A(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2b_1 _2056_ (.A_N(\scs.acc3_d2[2] ),
    .B(net358),
    .Y(_1723_));
 sky130_fd_sc_hd__a21oi_1 _2057_ (.A1(_1721_),
    .A2(_1723_),
    .B1(_1720_),
    .Y(_1724_));
 sky130_fd_sc_hd__a31o_1 _2058_ (.A1(_1720_),
    .A2(_1721_),
    .A3(_1723_),
    .B1(net80),
    .X(_1725_));
 sky130_fd_sc_hd__o221a_1 _2059_ (.A1(net668),
    .A2(net162),
    .B1(_1724_),
    .B2(_1725_),
    .C1(net483),
    .X(_0050_));
 sky130_fd_sc_hd__o21ai_1 _2060_ (.A1(_1720_),
    .A2(_1722_),
    .B1(_1723_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2b_1 _2061_ (.A_N(net357),
    .B(\scs.acc3_d2[3] ),
    .Y(_1727_));
 sky130_fd_sc_hd__inv_2 _2062_ (.A(_1727_),
    .Y(_1728_));
 sky130_fd_sc_hd__and2b_1 _2063_ (.A_N(\scs.acc3_d2[3] ),
    .B(net357),
    .X(_0315_));
 sky130_fd_sc_hd__o21a_1 _2064_ (.A1(_1728_),
    .A2(_0315_),
    .B1(_1726_),
    .X(_0316_));
 sky130_fd_sc_hd__o31ai_1 _2065_ (.A1(_1726_),
    .A2(_1728_),
    .A3(_0315_),
    .B1(net162),
    .Y(_0317_));
 sky130_fd_sc_hd__o221a_1 _2066_ (.A1(net678),
    .A2(net162),
    .B1(_0316_),
    .B2(_0317_),
    .C1(net488),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _2067_ (.A1(_1726_),
    .A2(_1727_),
    .B1(_0315_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_1 _2068_ (.A(net355),
    .B(\scs.acc3_d2[4] ),
    .Y(_0319_));
 sky130_fd_sc_hd__nand2_1 _2069_ (.A(_0318_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__or2_1 _2070_ (.A(_0318_),
    .B(_0319_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _2071_ (.A1(_0320_),
    .A2(_0321_),
    .B1(net82),
    .X(_0322_));
 sky130_fd_sc_hd__o211a_1 _2072_ (.A1(net702),
    .A2(net166),
    .B1(_0322_),
    .C1(net485),
    .X(_0052_));
 sky130_fd_sc_hd__nand2b_1 _2073_ (.A_N(net353),
    .B(\scs.acc3_d2[5] ),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2b_1 _2074_ (.A_N(\scs.acc3_d2[5] ),
    .B(net353),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _2075_ (.A(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _2076_ (.A(_0323_),
    .B(_0324_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _2077_ (.A(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21bo_1 _2078_ (.A1(net355),
    .A2(_1477_),
    .B1_N(_0320_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_1 _2079_ (.A(_0326_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21o_1 _2080_ (.A1(_0326_),
    .A2(_0328_),
    .B1(net82),
    .X(_0330_));
 sky130_fd_sc_hd__o221a_1 _2081_ (.A1(net742),
    .A2(net166),
    .B1(_0329_),
    .B2(_0330_),
    .C1(net488),
    .X(_0053_));
 sky130_fd_sc_hd__a31o_1 _2082_ (.A1(net355),
    .A2(_1477_),
    .A3(_0323_),
    .B1(_0325_),
    .X(_0331_));
 sky130_fd_sc_hd__a31o_1 _2083_ (.A1(_0318_),
    .A2(_0319_),
    .A3(_0327_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _2084_ (.A(net351),
    .B(_1476_),
    .Y(_0333_));
 sky130_fd_sc_hd__and2_1 _2085_ (.A(net351),
    .B(_1476_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_1 _2086_ (.A(_0333_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _2087_ (.A(_0332_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__or2_1 _2088_ (.A(_0332_),
    .B(_0335_),
    .X(_0337_));
 sky130_fd_sc_hd__a21o_1 _2089_ (.A1(_0336_),
    .A2(_0337_),
    .B1(net83),
    .X(_0338_));
 sky130_fd_sc_hd__o211a_1 _2090_ (.A1(net704),
    .A2(net167),
    .B1(_0338_),
    .C1(net486),
    .X(_0054_));
 sky130_fd_sc_hd__and2b_1 _2091_ (.A_N(net349),
    .B(\scs.acc3_d2[7] ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2b_1 _2092_ (.A_N(net349),
    .B(\scs.acc3_d2[7] ),
    .Y(_0340_));
 sky130_fd_sc_hd__and2b_1 _2093_ (.A_N(\scs.acc3_d2[7] ),
    .B(net349),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _2094_ (.A(_0339_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__a21oi_1 _2095_ (.A1(_0332_),
    .A2(_0335_),
    .B1(_0334_),
    .Y(_0343_));
 sky130_fd_sc_hd__o21ai_1 _2096_ (.A1(_0342_),
    .A2(_0343_),
    .B1(net167),
    .Y(_0344_));
 sky130_fd_sc_hd__a21o_1 _2097_ (.A1(_0342_),
    .A2(_0343_),
    .B1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o211a_1 _2098_ (.A1(net640),
    .A2(net167),
    .B1(_0345_),
    .C1(net500),
    .X(_0055_));
 sky130_fd_sc_hd__and2b_1 _2099_ (.A_N(\scs.acc3_d2[8] ),
    .B(net347),
    .X(_0346_));
 sky130_fd_sc_hd__nand2b_1 _2100_ (.A_N(net347),
    .B(\scs.acc3_d2[8] ),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2b_1 _2101_ (.A_N(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__a31o_1 _2102_ (.A1(net351),
    .A2(_1476_),
    .A3(_0340_),
    .B1(_0341_),
    .X(_0349_));
 sky130_fd_sc_hd__a31o_1 _2103_ (.A1(_0332_),
    .A2(_0335_),
    .A3(_0342_),
    .B1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__xnor2_1 _2104_ (.A(_0348_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__or2_1 _2105_ (.A(net676),
    .B(net182),
    .X(_0352_));
 sky130_fd_sc_hd__o211a_1 _2106_ (.A1(net98),
    .A2(_0351_),
    .B1(_0352_),
    .C1(net500),
    .X(_0056_));
 sky130_fd_sc_hd__and2b_1 _2107_ (.A_N(net345),
    .B(\scs.acc3_d2[9] ),
    .X(_0353_));
 sky130_fd_sc_hd__nand2b_1 _2108_ (.A_N(net345),
    .B(\scs.acc3_d2[9] ),
    .Y(_0354_));
 sky130_fd_sc_hd__and2b_1 _2109_ (.A_N(\scs.acc3_d2[9] ),
    .B(net345),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_1 _2110_ (.A(_0353_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_1 _2111_ (.A1(_0347_),
    .A2(_0350_),
    .B1(_0346_),
    .Y(_0357_));
 sky130_fd_sc_hd__and2_1 _2112_ (.A(_0356_),
    .B(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__o21ai_1 _2113_ (.A1(_0356_),
    .A2(_0357_),
    .B1(net182),
    .Y(_0359_));
 sky130_fd_sc_hd__o221a_1 _2114_ (.A1(net670),
    .A2(net182),
    .B1(_0358_),
    .B2(_0359_),
    .C1(net500),
    .X(_0057_));
 sky130_fd_sc_hd__nand2b_1 _2115_ (.A_N(\scs.acc3_d2[10] ),
    .B(net343),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _2116_ (.A(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2b_1 _2117_ (.A_N(net343),
    .B(\scs.acc3_d2[10] ),
    .Y(_0362_));
 sky130_fd_sc_hd__a211o_1 _2118_ (.A1(_0347_),
    .A2(_0350_),
    .B1(_0355_),
    .C1(_0346_),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _2119_ (.A1(_0360_),
    .A2(_0362_),
    .B1(_0363_),
    .B2(_0354_),
    .X(_0364_));
 sky130_fd_sc_hd__nand4_1 _2120_ (.A(_0354_),
    .B(_0360_),
    .C(_0362_),
    .D(_0363_),
    .Y(_0365_));
 sky130_fd_sc_hd__and3_1 _2121_ (.A(net183),
    .B(_0364_),
    .C(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a21oi_1 _2122_ (.A1(net690),
    .A2(net98),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _2123_ (.A(net574),
    .B(_0367_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _2124_ (.A(net653),
    .B(net98),
    .Y(_0368_));
 sky130_fd_sc_hd__and2b_1 _2125_ (.A_N(\scs.acc3_d2[11] ),
    .B(net341),
    .X(_0369_));
 sky130_fd_sc_hd__and2b_1 _2126_ (.A_N(net341),
    .B(\scs.acc3_d2[11] ),
    .X(_0370_));
 sky130_fd_sc_hd__a31oi_2 _2127_ (.A1(_0354_),
    .A2(_0362_),
    .A3(_0363_),
    .B1(_0361_),
    .Y(_0371_));
 sky130_fd_sc_hd__or3_1 _2128_ (.A(_0369_),
    .B(_0370_),
    .C(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__o21a_1 _2129_ (.A1(_0369_),
    .A2(_0370_),
    .B1(_0371_),
    .X(_0373_));
 sky130_fd_sc_hd__or3b_1 _2130_ (.A(_0373_),
    .B(net99),
    .C_N(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__a21oi_1 _2131_ (.A1(_0368_),
    .A2(_0374_),
    .B1(net574),
    .Y(_0059_));
 sky130_fd_sc_hd__o21ba_1 _2132_ (.A1(_0370_),
    .A2(_0371_),
    .B1_N(_0369_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2b_1 _2133_ (.A_N(net339),
    .B(\scs.acc3_d2[12] ),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2b_1 _2134_ (.A_N(\scs.acc3_d2[12] ),
    .B(net339),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(_0376_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__or2_1 _2136_ (.A(_0375_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _2137_ (.A(_0375_),
    .B(_0378_),
    .Y(_0380_));
 sky130_fd_sc_hd__and2_1 _2138_ (.A(_0379_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__or2_1 _2139_ (.A(net716),
    .B(net186),
    .X(_0382_));
 sky130_fd_sc_hd__o211a_1 _2140_ (.A1(net102),
    .A2(_0381_),
    .B1(_0382_),
    .C1(net504),
    .X(_0060_));
 sky130_fd_sc_hd__and2b_1 _2141_ (.A_N(net337),
    .B(\scs.acc3_d2[13] ),
    .X(_0383_));
 sky130_fd_sc_hd__nand2b_1 _2142_ (.A_N(\scs.acc3_d2[13] ),
    .B(net337),
    .Y(_0384_));
 sky130_fd_sc_hd__and2b_1 _2143_ (.A_N(_0383_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__inv_2 _2144_ (.A(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _2145_ (.A1(_0377_),
    .A2(_0379_),
    .B1(_0385_),
    .Y(_0387_));
 sky130_fd_sc_hd__a31o_1 _2146_ (.A1(_0377_),
    .A2(_0379_),
    .A3(_0385_),
    .B1(net102),
    .X(_0388_));
 sky130_fd_sc_hd__o221a_1 _2147_ (.A1(net772),
    .A2(net186),
    .B1(_0387_),
    .B2(_0388_),
    .C1(net504),
    .X(_0061_));
 sky130_fd_sc_hd__nand2b_1 _2148_ (.A_N(net335),
    .B(\scs.acc3_d2[14] ),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2b_1 _2149_ (.A_N(\scs.acc3_d2[14] ),
    .B(net335),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_1 _2150_ (.A(_0389_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__or3b_1 _2151_ (.A(\scs.acc3_d2[12] ),
    .B(_0383_),
    .C_N(net339),
    .X(_0392_));
 sky130_fd_sc_hd__o311a_1 _2152_ (.A1(_0375_),
    .A2(_0378_),
    .A3(_0386_),
    .B1(_0392_),
    .C1(_0384_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _2153_ (.A(_0391_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _2154_ (.A(_0391_),
    .B(_0393_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _2155_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _2156_ (.A(net731),
    .B(net186),
    .Y(_0397_));
 sky130_fd_sc_hd__a211oi_1 _2157_ (.A1(net187),
    .A2(_0396_),
    .B1(_0397_),
    .C1(net593),
    .Y(_0062_));
 sky130_fd_sc_hd__xnor2_2 _2158_ (.A(net333),
    .B(\scs.acc3_d2[15] ),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _2159_ (.A(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__a21oi_1 _2160_ (.A1(_0390_),
    .A2(_0394_),
    .B1(_0398_),
    .Y(_0400_));
 sky130_fd_sc_hd__a31o_1 _2161_ (.A1(_0390_),
    .A2(_0394_),
    .A3(_0398_),
    .B1(net102),
    .X(_0401_));
 sky130_fd_sc_hd__o221a_1 _2162_ (.A1(net658),
    .A2(net187),
    .B1(_0400_),
    .B2(_0401_),
    .C1(net505),
    .X(_0063_));
 sky130_fd_sc_hd__nand2b_1 _2163_ (.A_N(net331),
    .B(\scs.acc3_d2[16] ),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2b_1 _2164_ (.A_N(\scs.acc3_d2[16] ),
    .B(net331),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _2165_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21oi_1 _2166_ (.A1(_1474_),
    .A2(\scs.acc3_d2[15] ),
    .B1(\scs.acc3_d2[14] ),
    .Y(_0405_));
 sky130_fd_sc_hd__o2bb2a_1 _2167_ (.A1_N(net335),
    .A2_N(_0405_),
    .B1(\scs.acc3_d2[15] ),
    .B2(_1474_),
    .X(_0406_));
 sky130_fd_sc_hd__o31a_2 _2168_ (.A1(_0391_),
    .A2(_0393_),
    .A3(_0399_),
    .B1(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__xor2_1 _2169_ (.A(_0404_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _2170_ (.A(net682),
    .B(net203),
    .X(_0409_));
 sky130_fd_sc_hd__o211a_1 _2171_ (.A1(net115),
    .A2(_0408_),
    .B1(_0409_),
    .C1(net531),
    .X(_0064_));
 sky130_fd_sc_hd__and2b_1 _2172_ (.A_N(\scs.acc3_d2[17] ),
    .B(net329),
    .X(_0410_));
 sky130_fd_sc_hd__nand2b_1 _2173_ (.A_N(\scs.acc3_d2[17] ),
    .B(net329),
    .Y(_0411_));
 sky130_fd_sc_hd__and2b_1 _2174_ (.A_N(net329),
    .B(\scs.acc3_d2[17] ),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _2175_ (.A(_0410_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21a_1 _2176_ (.A1(_0404_),
    .A2(_0407_),
    .B1(_0403_),
    .X(_0414_));
 sky130_fd_sc_hd__xnor2_1 _2177_ (.A(_0413_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__or2_1 _2178_ (.A(net808),
    .B(net203),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_1 _2179_ (.A1(net115),
    .A2(_0415_),
    .B1(_0416_),
    .C1(net531),
    .X(_0065_));
 sky130_fd_sc_hd__nand2b_1 _2180_ (.A_N(\scs.acc3_d2[18] ),
    .B(net327),
    .Y(_0417_));
 sky130_fd_sc_hd__xnor2_2 _2181_ (.A(net327),
    .B(\scs.acc3_d2[18] ),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_2 _2182_ (.A(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__a21o_1 _2183_ (.A1(_0411_),
    .A2(_0414_),
    .B1(_0412_),
    .X(_0420_));
 sky130_fd_sc_hd__or2_1 _2184_ (.A(_0419_),
    .B(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__xnor2_1 _2185_ (.A(_0418_),
    .B(_0420_),
    .Y(_0422_));
 sky130_fd_sc_hd__or2_1 _2186_ (.A(net781),
    .B(net204),
    .X(_0423_));
 sky130_fd_sc_hd__o211a_1 _2187_ (.A1(net116),
    .A2(_0422_),
    .B1(_0423_),
    .C1(net533),
    .X(_0066_));
 sky130_fd_sc_hd__xnor2_1 _2188_ (.A(net325),
    .B(\scs.acc3_d2[19] ),
    .Y(_0424_));
 sky130_fd_sc_hd__a21oi_1 _2189_ (.A1(_0417_),
    .A2(_0421_),
    .B1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a31o_1 _2190_ (.A1(_0417_),
    .A2(_0421_),
    .A3(_0424_),
    .B1(net118),
    .X(_0426_));
 sky130_fd_sc_hd__o221a_1 _2191_ (.A1(net652),
    .A2(net204),
    .B1(_0425_),
    .B2(_0426_),
    .C1(net531),
    .X(_0067_));
 sky130_fd_sc_hd__and2b_1 _2192_ (.A_N(net323),
    .B(\scs.acc3_d2[20] ),
    .X(_0427_));
 sky130_fd_sc_hd__and2b_1 _2193_ (.A_N(\scs.acc3_d2[20] ),
    .B(net323),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _2194_ (.A(_0427_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _2195_ (.A(_0418_),
    .B(_0424_),
    .Y(_0430_));
 sky130_fd_sc_hd__a211o_1 _2196_ (.A1(_0403_),
    .A2(_0411_),
    .B1(_0412_),
    .C1(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__a21o_1 _2197_ (.A1(_1473_),
    .A2(\scs.acc3_d2[19] ),
    .B1(_0417_),
    .X(_0432_));
 sky130_fd_sc_hd__o211a_1 _2198_ (.A1(_1473_),
    .A2(\scs.acc3_d2[19] ),
    .B1(_0431_),
    .C1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__or4_1 _2199_ (.A(_0404_),
    .B(_0410_),
    .C(_0412_),
    .D(_0430_),
    .X(_0434_));
 sky130_fd_sc_hd__o21ai_1 _2200_ (.A1(_0407_),
    .A2(_0434_),
    .B1(_0433_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _2201_ (.A(_0429_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _2202_ (.A(net665),
    .B(net208),
    .Y(_0437_));
 sky130_fd_sc_hd__a211oi_1 _2203_ (.A1(net208),
    .A2(_0436_),
    .B1(_0437_),
    .C1(net593),
    .Y(_0068_));
 sky130_fd_sc_hd__and2b_1 _2204_ (.A_N(\scs.acc3_d2[21] ),
    .B(net321),
    .X(_0438_));
 sky130_fd_sc_hd__nand2b_1 _2205_ (.A_N(\scs.acc3_d2[21] ),
    .B(net321),
    .Y(_0439_));
 sky130_fd_sc_hd__and2b_1 _2206_ (.A_N(net321),
    .B(\scs.acc3_d2[21] ),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _2207_ (.A(_0438_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a21oi_1 _2208_ (.A1(_0429_),
    .A2(_0435_),
    .B1(_0428_),
    .Y(_0442_));
 sky130_fd_sc_hd__and2_1 _2209_ (.A(_0441_),
    .B(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__o21ai_1 _2210_ (.A1(_0441_),
    .A2(_0442_),
    .B1(net210),
    .Y(_0444_));
 sky130_fd_sc_hd__o221a_1 _2211_ (.A1(net654),
    .A2(net207),
    .B1(_0443_),
    .B2(_0444_),
    .C1(net533),
    .X(_0069_));
 sky130_fd_sc_hd__nand2b_1 _2212_ (.A_N(net319),
    .B(\scs.acc3_d2[22] ),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2b_1 _2213_ (.A_N(\scs.acc3_d2[22] ),
    .B(net319),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _2214_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__a21o_1 _2215_ (.A1(_0439_),
    .A2(_0442_),
    .B1(_0440_),
    .X(_0448_));
 sky130_fd_sc_hd__xnor2_1 _2216_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(net207),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__o211a_1 _2218_ (.A1(net753),
    .A2(net223),
    .B1(_0450_),
    .C1(net547),
    .X(_0070_));
 sky130_fd_sc_hd__and2b_1 _2219_ (.A_N(net318),
    .B(\scs.acc3_d2[23] ),
    .X(_0451_));
 sky130_fd_sc_hd__and2b_1 _2220_ (.A_N(\scs.acc3_d2[23] ),
    .B(net318),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_1 _2221_ (.A1(_0447_),
    .A2(_0448_),
    .B1(_0446_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21ai_1 _2222_ (.A1(_0451_),
    .A2(_0452_),
    .B1(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o31a_1 _2223_ (.A1(_0451_),
    .A2(_0452_),
    .A3(_0453_),
    .B1(net210),
    .X(_0455_));
 sky130_fd_sc_hd__a221oi_1 _2224_ (.A1(_1463_),
    .A2(net119),
    .B1(_0454_),
    .B2(_0455_),
    .C1(net607),
    .Y(_0071_));
 sky130_fd_sc_hd__nand2b_1 _2225_ (.A_N(\scs.acc3_d2[24] ),
    .B(net316),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2b_1 _2226_ (.A_N(net316),
    .B(\scs.acc3_d2[24] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _2227_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__or3_1 _2228_ (.A(_0447_),
    .B(_0451_),
    .C(_0452_),
    .X(_0459_));
 sky130_fd_sc_hd__or4b_1 _2229_ (.A(_0438_),
    .B(_0440_),
    .C(_0459_),
    .D_N(_0429_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2b_1 _2230_ (.A_N(_0440_),
    .B(_0428_),
    .Y(_0461_));
 sky130_fd_sc_hd__a21o_1 _2231_ (.A1(_0439_),
    .A2(_0461_),
    .B1(_0459_),
    .X(_0462_));
 sky130_fd_sc_hd__o21ba_1 _2232_ (.A1(_0446_),
    .A2(_0451_),
    .B1_N(_0452_),
    .X(_0463_));
 sky130_fd_sc_hd__o211a_1 _2233_ (.A1(_0433_),
    .A2(_0460_),
    .B1(_0462_),
    .C1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__o31a_1 _2234_ (.A1(_0407_),
    .A2(_0434_),
    .A3(_0460_),
    .B1(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__or2_1 _2235_ (.A(_0458_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_1 _2236_ (.A(_0458_),
    .B(_0465_),
    .Y(_0467_));
 sky130_fd_sc_hd__and2_1 _2237_ (.A(_0466_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__or2_1 _2238_ (.A(net686),
    .B(net223),
    .X(_0469_));
 sky130_fd_sc_hd__o211a_1 _2239_ (.A1(net134),
    .A2(_0468_),
    .B1(_0469_),
    .C1(net549),
    .X(_0072_));
 sky130_fd_sc_hd__nand2b_1 _2240_ (.A_N(\scs.acc3_d2[25] ),
    .B(net315),
    .Y(_0470_));
 sky130_fd_sc_hd__and2b_1 _2241_ (.A_N(net315),
    .B(\scs.acc3_d2[25] ),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _2242_ (.A(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _2243_ (.A(_0470_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__and2_1 _2244_ (.A(_0456_),
    .B(_0466_),
    .X(_0474_));
 sky130_fd_sc_hd__xor2_1 _2245_ (.A(_0473_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__or2_1 _2246_ (.A(net688),
    .B(net224),
    .X(_0476_));
 sky130_fd_sc_hd__o211a_1 _2247_ (.A1(net135),
    .A2(_0475_),
    .B1(_0476_),
    .C1(net547),
    .X(_0073_));
 sky130_fd_sc_hd__nand2b_1 _2248_ (.A_N(\scs.acc3_d2[26] ),
    .B(net313),
    .Y(_0477_));
 sky130_fd_sc_hd__xnor2_2 _2249_ (.A(net313),
    .B(\scs.acc3_d2[26] ),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _2250_ (.A(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a31o_1 _2251_ (.A1(_0456_),
    .A2(_0466_),
    .A3(_0470_),
    .B1(_0471_),
    .X(_0480_));
 sky130_fd_sc_hd__or2_1 _2252_ (.A(_0479_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_1 _2253_ (.A(_0478_),
    .B(_0480_),
    .Y(_0482_));
 sky130_fd_sc_hd__or2_1 _2254_ (.A(\scs.diff1[26] ),
    .B(net227),
    .X(_0483_));
 sky130_fd_sc_hd__o211a_1 _2255_ (.A1(net139),
    .A2(_0482_),
    .B1(_0483_),
    .C1(net552),
    .X(_0074_));
 sky130_fd_sc_hd__xnor2_1 _2256_ (.A(net311),
    .B(\scs.acc3_d2[27] ),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _2257_ (.A1(_0477_),
    .A2(_0481_),
    .B1(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__a31o_1 _2258_ (.A1(_0477_),
    .A2(_0481_),
    .A3(_0484_),
    .B1(net136),
    .X(_0486_));
 sky130_fd_sc_hd__o221a_1 _2259_ (.A1(net854),
    .A2(net227),
    .B1(_0485_),
    .B2(_0486_),
    .C1(net547),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _2260_ (.A(_0478_),
    .B(_0484_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21o_1 _2261_ (.A1(_0456_),
    .A2(_0470_),
    .B1(_0471_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_1 _2262_ (.A1(_1472_),
    .A2(\scs.acc3_d2[27] ),
    .B1(_0477_),
    .X(_0489_));
 sky130_fd_sc_hd__o221a_1 _2263_ (.A1(_1472_),
    .A2(\scs.acc3_d2[27] ),
    .B1(_0487_),
    .B2(_0488_),
    .C1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__o31a_1 _2264_ (.A1(_0466_),
    .A2(_0473_),
    .A3(_0487_),
    .B1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__and2b_1 _2265_ (.A_N(net310),
    .B(\scs.acc3_d2[28] ),
    .X(_0492_));
 sky130_fd_sc_hd__nand2b_1 _2266_ (.A_N(\scs.acc3_d2[28] ),
    .B(net310),
    .Y(_0493_));
 sky130_fd_sc_hd__and2b_1 _2267_ (.A_N(_0492_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _2268_ (.A(_0491_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__o21ai_1 _2269_ (.A1(_0491_),
    .A2(_0494_),
    .B1(net229),
    .Y(_0496_));
 sky130_fd_sc_hd__o221a_1 _2270_ (.A1(net765),
    .A2(net227),
    .B1(_0495_),
    .B2(_0496_),
    .C1(net552),
    .X(_0076_));
 sky130_fd_sc_hd__o21ai_1 _2271_ (.A1(_0491_),
    .A2(_0492_),
    .B1(_0493_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2b_1 _2272_ (.A_N(net309),
    .B(\scs.acc3_d2[29] ),
    .Y(_0498_));
 sky130_fd_sc_hd__and2b_1 _2273_ (.A_N(\scs.acc3_d2[29] ),
    .B(net309),
    .X(_0499_));
 sky130_fd_sc_hd__inv_2 _2274_ (.A(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _2275_ (.A(_0498_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_1 _2276_ (.A(_0497_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21o_1 _2277_ (.A1(_0497_),
    .A2(_0501_),
    .B1(net141),
    .X(_0503_));
 sky130_fd_sc_hd__o221a_1 _2278_ (.A1(net726),
    .A2(net230),
    .B1(_0502_),
    .B2(_0503_),
    .C1(net552),
    .X(_0077_));
 sky130_fd_sc_hd__nand2b_1 _2279_ (.A_N(\scs.acc3_d2[30] ),
    .B(net695),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2b_1 _2280_ (.A_N(net695),
    .B(\scs.acc3_d2[30] ),
    .Y(_0505_));
 sky130_fd_sc_hd__a21o_1 _2281_ (.A1(_0497_),
    .A2(_0498_),
    .B1(_0499_),
    .X(_0506_));
 sky130_fd_sc_hd__a21o_1 _2282_ (.A1(_0504_),
    .A2(_0505_),
    .B1(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a31oi_1 _2283_ (.A1(_0504_),
    .A2(_0505_),
    .A3(_0506_),
    .B1(net142),
    .Y(_0508_));
 sky130_fd_sc_hd__a22o_1 _2284_ (.A1(net720),
    .A2(net141),
    .B1(_0507_),
    .B2(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _2285_ (.A(net553),
    .B(_0509_),
    .X(_0078_));
 sky130_fd_sc_hd__a21bo_1 _2286_ (.A1(_0505_),
    .A2(_0506_),
    .B1_N(_0504_),
    .X(_0510_));
 sky130_fd_sc_hd__xor2_1 _2287_ (.A(\scs.acc3[31] ),
    .B(\scs.acc3_d2[31] ),
    .X(_0511_));
 sky130_fd_sc_hd__xnor2_1 _2288_ (.A(_0510_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__or2_1 _2289_ (.A(net661),
    .B(net230),
    .X(_0513_));
 sky130_fd_sc_hd__o211a_1 _2290_ (.A1(net141),
    .A2(_0512_),
    .B1(_0513_),
    .C1(net553),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _2291_ (.A(net789),
    .B(net163),
    .X(_0514_));
 sky130_fd_sc_hd__o211a_1 _2292_ (.A1(net806),
    .A2(net80),
    .B1(_0514_),
    .C1(net483),
    .X(_0080_));
 sky130_fd_sc_hd__or2_1 _2293_ (.A(net801),
    .B(net163),
    .X(_0515_));
 sky130_fd_sc_hd__o211a_1 _2294_ (.A1(net359),
    .A2(net80),
    .B1(_0515_),
    .C1(net483),
    .X(_0081_));
 sky130_fd_sc_hd__or2_1 _2295_ (.A(net782),
    .B(net164),
    .X(_0516_));
 sky130_fd_sc_hd__o211a_1 _2296_ (.A1(net358),
    .A2(net80),
    .B1(_0516_),
    .C1(net510),
    .X(_0082_));
 sky130_fd_sc_hd__or2_1 _2297_ (.A(net787),
    .B(net164),
    .X(_0517_));
 sky130_fd_sc_hd__o211a_1 _2298_ (.A1(net357),
    .A2(net86),
    .B1(_0517_),
    .C1(net487),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_1 _2299_ (.A(_1477_),
    .B(net84),
    .Y(_0518_));
 sky130_fd_sc_hd__o211a_1 _2300_ (.A1(net355),
    .A2(net84),
    .B1(_0518_),
    .C1(net487),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _2301_ (.A(net788),
    .B(net169),
    .X(_0519_));
 sky130_fd_sc_hd__o211a_1 _2302_ (.A1(net353),
    .A2(net84),
    .B1(_0519_),
    .C1(net509),
    .X(_0085_));
 sky130_fd_sc_hd__or2_1 _2303_ (.A(net709),
    .B(net168),
    .X(_0520_));
 sky130_fd_sc_hd__o211a_1 _2304_ (.A1(net351),
    .A2(net85),
    .B1(_0520_),
    .C1(net502),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _2305_ (.A(net834),
    .B(net168),
    .X(_0521_));
 sky130_fd_sc_hd__o211a_1 _2306_ (.A1(net349),
    .A2(net84),
    .B1(_0521_),
    .C1(net502),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _2307_ (.A(net760),
    .B(net184),
    .X(_0522_));
 sky130_fd_sc_hd__o211a_1 _2308_ (.A1(net347),
    .A2(net100),
    .B1(_0522_),
    .C1(net503),
    .X(_0088_));
 sky130_fd_sc_hd__or2_1 _2309_ (.A(net821),
    .B(net184),
    .X(_0523_));
 sky130_fd_sc_hd__o211a_1 _2310_ (.A1(net345),
    .A2(net100),
    .B1(_0523_),
    .C1(net502),
    .X(_0089_));
 sky130_fd_sc_hd__or2_1 _2311_ (.A(net799),
    .B(net185),
    .X(_0524_));
 sky130_fd_sc_hd__o211a_1 _2312_ (.A1(net343),
    .A2(net101),
    .B1(_0524_),
    .C1(net502),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _2313_ (.A(net795),
    .B(net185),
    .X(_0525_));
 sky130_fd_sc_hd__o211a_1 _2314_ (.A1(net341),
    .A2(net101),
    .B1(_0525_),
    .C1(net505),
    .X(_0091_));
 sky130_fd_sc_hd__or2_1 _2315_ (.A(net790),
    .B(net188),
    .X(_0526_));
 sky130_fd_sc_hd__o211a_1 _2316_ (.A1(net339),
    .A2(net104),
    .B1(_0526_),
    .C1(net505),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _2317_ (.A(net791),
    .B(net188),
    .X(_0527_));
 sky130_fd_sc_hd__o211a_1 _2318_ (.A1(net337),
    .A2(net104),
    .B1(_0527_),
    .C1(net505),
    .X(_0093_));
 sky130_fd_sc_hd__or2_1 _2319_ (.A(net761),
    .B(net189),
    .X(_0528_));
 sky130_fd_sc_hd__o211a_1 _2320_ (.A1(net335),
    .A2(net103),
    .B1(_0528_),
    .C1(net531),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _2321_ (.A(net858),
    .B(net189),
    .X(_0529_));
 sky130_fd_sc_hd__o211a_1 _2322_ (.A1(net333),
    .A2(net103),
    .B1(_0529_),
    .C1(net558),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _2323_ (.A(net810),
    .B(net205),
    .X(_0530_));
 sky130_fd_sc_hd__o211a_1 _2324_ (.A1(net331),
    .A2(net117),
    .B1(_0530_),
    .C1(net558),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _2325_ (.A(net811),
    .B(net205),
    .X(_0531_));
 sky130_fd_sc_hd__o211a_1 _2326_ (.A1(net329),
    .A2(net117),
    .B1(_0531_),
    .C1(net560),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _2327_ (.A(net859),
    .B(net206),
    .X(_0532_));
 sky130_fd_sc_hd__o211a_1 _2328_ (.A1(net327),
    .A2(net117),
    .B1(_0532_),
    .C1(net561),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _2329_ (.A(net864),
    .B(net206),
    .X(_0533_));
 sky130_fd_sc_hd__o211a_1 _2330_ (.A1(net325),
    .A2(net117),
    .B1(_0533_),
    .C1(net533),
    .X(_0099_));
 sky130_fd_sc_hd__or2_1 _2331_ (.A(net771),
    .B(net209),
    .X(_0534_));
 sky130_fd_sc_hd__o211a_1 _2332_ (.A1(net323),
    .A2(net119),
    .B1(_0534_),
    .C1(net561),
    .X(_0100_));
 sky130_fd_sc_hd__or2_1 _2333_ (.A(net819),
    .B(net209),
    .X(_0535_));
 sky130_fd_sc_hd__o211a_1 _2334_ (.A1(net321),
    .A2(net120),
    .B1(_0535_),
    .C1(net533),
    .X(_0101_));
 sky130_fd_sc_hd__or2_1 _2335_ (.A(net755),
    .B(net209),
    .X(_0536_));
 sky130_fd_sc_hd__o211a_1 _2336_ (.A1(net319),
    .A2(net120),
    .B1(_0536_),
    .C1(net564),
    .X(_0102_));
 sky130_fd_sc_hd__or2_1 _2337_ (.A(net798),
    .B(net209),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _2338_ (.A1(net318),
    .A2(net120),
    .B1(_0537_),
    .C1(net564),
    .X(_0103_));
 sky130_fd_sc_hd__or2_1 _2339_ (.A(net797),
    .B(net225),
    .X(_0538_));
 sky130_fd_sc_hd__o211a_1 _2340_ (.A1(net316),
    .A2(net137),
    .B1(_0538_),
    .C1(net547),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _2341_ (.A(net779),
    .B(net225),
    .X(_0539_));
 sky130_fd_sc_hd__o211a_1 _2342_ (.A1(net315),
    .A2(net137),
    .B1(_0539_),
    .C1(net564),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _2343_ (.A(net861),
    .B(net226),
    .X(_0540_));
 sky130_fd_sc_hd__o211a_1 _2344_ (.A1(net313),
    .A2(net143),
    .B1(_0540_),
    .C1(net567),
    .X(_0106_));
 sky130_fd_sc_hd__or2_1 _2345_ (.A(net862),
    .B(net226),
    .X(_0541_));
 sky130_fd_sc_hd__o211a_1 _2346_ (.A1(net311),
    .A2(net136),
    .B1(_0541_),
    .C1(net565),
    .X(_0107_));
 sky130_fd_sc_hd__or2_1 _2347_ (.A(net780),
    .B(net229),
    .X(_0542_));
 sky130_fd_sc_hd__o211a_1 _2348_ (.A1(net310),
    .A2(net143),
    .B1(_0542_),
    .C1(net552),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _2349_ (.A(net774),
    .B(net229),
    .X(_0543_));
 sky130_fd_sc_hd__o211a_1 _2350_ (.A1(net309),
    .A2(net143),
    .B1(_0543_),
    .C1(net567),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _2351_ (.A(net796),
    .B(net229),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _2352_ (.A1(net792),
    .A2(net142),
    .B1(_0544_),
    .C1(net567),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _2353_ (.A(net793),
    .B(net230),
    .X(_0545_));
 sky130_fd_sc_hd__o211a_1 _2354_ (.A1(\scs.acc3[31] ),
    .A2(net141),
    .B1(_0545_),
    .C1(net567),
    .X(_0111_));
 sky130_fd_sc_hd__o22a_1 _2355_ (.A1(_1455_),
    .A2(\scs.oversample_in[1] ),
    .B1(\scs.oversample_in[5] ),
    .B2(_1451_),
    .X(_0546_));
 sky130_fd_sc_hd__o221a_1 _2356_ (.A1(net270),
    .A2(_1479_),
    .B1(\scs.oversample_in[2] ),
    .B2(_1454_),
    .C1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o21ai_1 _2357_ (.A1(_1452_),
    .A2(\scs.oversample_in[4] ),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a221o_1 _2358_ (.A1(net260),
    .A2(_1482_),
    .B1(_1483_),
    .B2(net256),
    .C1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__o22a_1 _2359_ (.A1(_1453_),
    .A2(\scs.oversample_in[3] ),
    .B1(_1483_),
    .B2(net256),
    .X(_0550_));
 sky130_fd_sc_hd__o21ai_1 _2360_ (.A1(net260),
    .A2(_1482_),
    .B1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__a22o_1 _2361_ (.A1(_1452_),
    .A2(\scs.oversample_in[4] ),
    .B1(\scs.oversample_in[5] ),
    .B2(_1451_),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _2362_ (.A1(_1454_),
    .A2(\scs.oversample_in[2] ),
    .B1(\scs.oversample_in[9] ),
    .B2(_1449_),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _2363_ (.A1(_1450_),
    .A2(\scs.oversample_in[7] ),
    .B1(_1484_),
    .B2(\scs.word_count[8] ),
    .X(_0554_));
 sky130_fd_sc_hd__o22a_1 _2364_ (.A1(net267),
    .A2(_1481_),
    .B1(\scs.oversample_in[7] ),
    .B2(_1450_),
    .X(_0555_));
 sky130_fd_sc_hd__or4b_1 _2365_ (.A(_0552_),
    .B(_0553_),
    .C(_0554_),
    .D_N(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__or4_1 _2366_ (.A(net254),
    .B(_0549_),
    .C(_0551_),
    .D(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_1 _2367_ (.A(net427),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__o211a_1 _2368_ (.A1(net427),
    .A2(net636),
    .B1(net509),
    .C1(_0558_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _2369_ (.A(\scs.acc1[0] ),
    .B(net412),
    .X(_0559_));
 sky130_fd_sc_hd__a21oi_1 _2370_ (.A1(net436),
    .A2(\scs.acc1[0] ),
    .B1(net637),
    .Y(_0560_));
 sky130_fd_sc_hd__a211oi_1 _2371_ (.A1(net436),
    .A2(net880),
    .B1(net638),
    .C1(net582),
    .Y(_0113_));
 sky130_fd_sc_hd__nand2_1 _2372_ (.A(net308),
    .B(net411),
    .Y(_0561_));
 sky130_fd_sc_hd__or2_1 _2373_ (.A(net308),
    .B(net411),
    .X(_0562_));
 sky130_fd_sc_hd__and3_1 _2374_ (.A(_0559_),
    .B(_0561_),
    .C(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a21oi_1 _2375_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0559_),
    .Y(_0564_));
 sky130_fd_sc_hd__o21ai_1 _2376_ (.A1(_0563_),
    .A2(_0564_),
    .B1(net437),
    .Y(_0565_));
 sky130_fd_sc_hd__o211a_1 _2377_ (.A1(net436),
    .A2(net624),
    .B1(net514),
    .C1(_0565_),
    .X(_0114_));
 sky130_fd_sc_hd__a21boi_2 _2378_ (.A1(_0559_),
    .A2(_0562_),
    .B1_N(_0561_),
    .Y(_0566_));
 sky130_fd_sc_hd__nor2_1 _2379_ (.A(net306),
    .B(net409),
    .Y(_0567_));
 sky130_fd_sc_hd__or2_1 _2380_ (.A(net306),
    .B(net410),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _2381_ (.A(net306),
    .B(net410),
    .Y(_0569_));
 sky130_fd_sc_hd__a21oi_1 _2382_ (.A1(_0568_),
    .A2(_0569_),
    .B1(_0566_),
    .Y(_0570_));
 sky130_fd_sc_hd__a31o_1 _2383_ (.A1(_0566_),
    .A2(_0568_),
    .A3(_0569_),
    .B1(net241),
    .X(_0571_));
 sky130_fd_sc_hd__nor2_1 _2384_ (.A(net434),
    .B(net409),
    .Y(_0572_));
 sky130_fd_sc_hd__o221a_1 _2385_ (.A1(net436),
    .A2(net872),
    .B1(_0570_),
    .B2(_0571_),
    .C1(net514),
    .X(_0115_));
 sky130_fd_sc_hd__o21a_1 _2386_ (.A1(_0566_),
    .A2(_0567_),
    .B1(_0569_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_1 _2387_ (.A(net304),
    .B(net407),
    .Y(_0574_));
 sky130_fd_sc_hd__or2_1 _2388_ (.A(net304),
    .B(net408),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _2389_ (.A(net304),
    .B(net408),
    .Y(_0576_));
 sky130_fd_sc_hd__a21oi_1 _2390_ (.A1(_0575_),
    .A2(_0576_),
    .B1(_0573_),
    .Y(_0577_));
 sky130_fd_sc_hd__a31o_1 _2391_ (.A1(_0573_),
    .A2(_0575_),
    .A3(_0576_),
    .B1(net241),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_1 _2392_ (.A(net438),
    .B(net407),
    .Y(_0579_));
 sky130_fd_sc_hd__o221a_1 _2393_ (.A1(net438),
    .A2(net870),
    .B1(_0577_),
    .B2(_0578_),
    .C1(net514),
    .X(_0116_));
 sky130_fd_sc_hd__o21ai_2 _2394_ (.A1(_0573_),
    .A2(_0574_),
    .B1(_0576_),
    .Y(_0580_));
 sky130_fd_sc_hd__and2_1 _2395_ (.A(net303),
    .B(net405),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _2396_ (.A(net303),
    .B(net406),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _2397_ (.A(_0581_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__xor2_1 _2398_ (.A(net609),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _2399_ (.A(net431),
    .B(net406),
    .X(_0585_));
 sky130_fd_sc_hd__o211a_1 _2400_ (.A1(net237),
    .A2(_0584_),
    .B1(_0585_),
    .C1(net509),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _2401_ (.A(net300),
    .B(net404),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _2402_ (.A(net300),
    .B(net404),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_2 _2403_ (.A(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__and2_1 _2404_ (.A(_0586_),
    .B(_0587_),
    .X(_0589_));
 sky130_fd_sc_hd__a21oi_1 _2405_ (.A1(_0580_),
    .A2(_0583_),
    .B1(_0581_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _2406_ (.A(_0589_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o21a_1 _2407_ (.A1(_0589_),
    .A2(_0590_),
    .B1(net431),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _2408_ (.A(net431),
    .B(net403),
    .Y(_0593_));
 sky130_fd_sc_hd__a211oi_1 _2409_ (.A1(_0591_),
    .A2(_0592_),
    .B1(_0593_),
    .C1(net578),
    .Y(_0118_));
 sky130_fd_sc_hd__a31o_1 _2410_ (.A1(net303),
    .A2(net406),
    .A3(_0586_),
    .B1(_0588_),
    .X(_0594_));
 sky130_fd_sc_hd__a31o_4 _2411_ (.A1(_0580_),
    .A2(_0583_),
    .A3(_0589_),
    .B1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _2412_ (.A(net298),
    .B(net401),
    .Y(_0596_));
 sky130_fd_sc_hd__or2_1 _2413_ (.A(net298),
    .B(net402),
    .X(_0597_));
 sky130_fd_sc_hd__nand2_1 _2414_ (.A(_0596_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _2415_ (.A(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__xnor2_1 _2416_ (.A(_0595_),
    .B(_0598_),
    .Y(_0600_));
 sky130_fd_sc_hd__or2_1 _2417_ (.A(net432),
    .B(net402),
    .X(_0601_));
 sky130_fd_sc_hd__o211a_1 _2418_ (.A1(net236),
    .A2(_0600_),
    .B1(_0601_),
    .C1(net517),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _2419_ (.A(\scs.acc1[7] ),
    .B(net400),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_1 _2420_ (.A(\scs.acc1[7] ),
    .B(net400),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _2421_ (.A(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__and2_1 _2422_ (.A(_0602_),
    .B(_0603_),
    .X(_0605_));
 sky130_fd_sc_hd__a21boi_1 _2423_ (.A1(_0595_),
    .A2(_0599_),
    .B1_N(_0596_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _2424_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__o21a_1 _2425_ (.A1(_0605_),
    .A2(_0606_),
    .B1(net431),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _2426_ (.A(net430),
    .B(net399),
    .Y(_0609_));
 sky130_fd_sc_hd__a211oi_1 _2427_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0609_),
    .C1(net586),
    .Y(_0120_));
 sky130_fd_sc_hd__a31o_1 _2428_ (.A1(net298),
    .A2(net402),
    .A3(_0602_),
    .B1(_0604_),
    .X(_0610_));
 sky130_fd_sc_hd__a31oi_4 _2429_ (.A1(_0595_),
    .A2(_0599_),
    .A3(_0605_),
    .B1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand2_1 _2430_ (.A(net297),
    .B(net397),
    .Y(_0612_));
 sky130_fd_sc_hd__or2_1 _2431_ (.A(net297),
    .B(net398),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(_0612_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__xor2_1 _2433_ (.A(_0611_),
    .B(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or2_1 _2434_ (.A(net442),
    .B(net398),
    .X(_0616_));
 sky130_fd_sc_hd__o211a_1 _2435_ (.A1(net243),
    .A2(_0615_),
    .B1(_0616_),
    .C1(net516),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _2436_ (.A(net294),
    .B(net395),
    .Y(_0617_));
 sky130_fd_sc_hd__and2_1 _2437_ (.A(net294),
    .B(net396),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _2438_ (.A(net294),
    .B(net396),
    .Y(_0619_));
 sky130_fd_sc_hd__o21ai_1 _2439_ (.A1(_0611_),
    .A2(_0614_),
    .B1(_0612_),
    .Y(_0620_));
 sky130_fd_sc_hd__o21ai_1 _2440_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__o31a_1 _2441_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0620_),
    .B1(net442),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _2442_ (.A(net441),
    .B(net395),
    .Y(_0623_));
 sky130_fd_sc_hd__a211oi_1 _2443_ (.A1(_0621_),
    .A2(_0622_),
    .B1(_0623_),
    .C1(net586),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(net293),
    .B(\scs.acc2[10] ),
    .Y(_0624_));
 sky130_fd_sc_hd__or2_1 _2445_ (.A(net293),
    .B(net394),
    .X(_0625_));
 sky130_fd_sc_hd__inv_2 _2446_ (.A(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _2447_ (.A(_0624_),
    .B(_0625_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand3b_1 _2448_ (.A_N(_0617_),
    .B(net398),
    .C(net297),
    .Y(_0628_));
 sky130_fd_sc_hd__o311a_4 _2449_ (.A1(_0611_),
    .A2(_0614_),
    .A3(_0617_),
    .B1(_0619_),
    .C1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__xor2_1 _2450_ (.A(_0627_),
    .B(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(net394),
    .A1(_0630_),
    .S(net442),
    .X(_0631_));
 sky130_fd_sc_hd__and2_1 _2452_ (.A(net516),
    .B(_0631_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_1 _2453_ (.A(\scs.acc1[11] ),
    .B(net393),
    .Y(_0632_));
 sky130_fd_sc_hd__or2_1 _2454_ (.A(\scs.acc1[11] ),
    .B(net393),
    .X(_0633_));
 sky130_fd_sc_hd__and2_1 _2455_ (.A(_0632_),
    .B(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__o21ai_4 _2456_ (.A1(_0626_),
    .A2(_0629_),
    .B1(_0624_),
    .Y(_0635_));
 sky130_fd_sc_hd__o21ai_1 _2457_ (.A1(_0634_),
    .A2(_0635_),
    .B1(net445),
    .Y(_0636_));
 sky130_fd_sc_hd__a21oi_1 _2458_ (.A1(_0634_),
    .A2(_0635_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _2459_ (.A1(net243),
    .A2(net629),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _2460_ (.A(net587),
    .B(_0638_),
    .Y(_0124_));
 sky130_fd_sc_hd__a21boi_2 _2461_ (.A1(_0633_),
    .A2(_0635_),
    .B1_N(_0632_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _2462_ (.A(net291),
    .B(net391),
    .Y(_0640_));
 sky130_fd_sc_hd__or2_1 _2463_ (.A(net291),
    .B(net392),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_1 _2464_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__xor2_1 _2465_ (.A(_0639_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__or2_1 _2466_ (.A(net445),
    .B(net392),
    .X(_0644_));
 sky130_fd_sc_hd__o211a_1 _2467_ (.A1(net244),
    .A2(_0643_),
    .B1(_0644_),
    .C1(net517),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _2468_ (.A(net290),
    .B(net390),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_1 _2469_ (.A(net290),
    .B(net390),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _2470_ (.A(_0645_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__o21ai_1 _2471_ (.A1(_0639_),
    .A2(_0642_),
    .B1(_0640_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _2472_ (.A(_0647_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__o21a_1 _2473_ (.A1(_0647_),
    .A2(_0648_),
    .B1(net445),
    .X(_0650_));
 sky130_fd_sc_hd__nor2_1 _2474_ (.A(net443),
    .B(net389),
    .Y(_0651_));
 sky130_fd_sc_hd__a211oi_1 _2475_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0651_),
    .C1(net587),
    .Y(_0126_));
 sky130_fd_sc_hd__and2_1 _2476_ (.A(net287),
    .B(net387),
    .X(_0652_));
 sky130_fd_sc_hd__nor2_1 _2477_ (.A(net287),
    .B(net388),
    .Y(_0653_));
 sky130_fd_sc_hd__or2_1 _2478_ (.A(_0652_),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nand3_1 _2479_ (.A(net291),
    .B(net392),
    .C(_0645_),
    .Y(_0655_));
 sky130_fd_sc_hd__o311a_4 _2480_ (.A1(_0639_),
    .A2(_0642_),
    .A3(_0647_),
    .B1(_0655_),
    .C1(_0646_),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _2481_ (.A(_0654_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__xor2_1 _2482_ (.A(_0654_),
    .B(_0656_),
    .X(_0658_));
 sky130_fd_sc_hd__or2_1 _2483_ (.A(net446),
    .B(net388),
    .X(_0659_));
 sky130_fd_sc_hd__o211a_1 _2484_ (.A1(net244),
    .A2(_0658_),
    .B1(_0659_),
    .C1(net559),
    .X(_0127_));
 sky130_fd_sc_hd__xnor2_1 _2485_ (.A(net283),
    .B(net386),
    .Y(_0660_));
 sky130_fd_sc_hd__or3_1 _2486_ (.A(_0652_),
    .B(_0657_),
    .C(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__o21ai_1 _2487_ (.A1(_0652_),
    .A2(_0657_),
    .B1(_0660_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_1 _2488_ (.A(net446),
    .B(net385),
    .Y(_0663_));
 sky130_fd_sc_hd__a311oi_1 _2489_ (.A1(net445),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0663_),
    .C1(net594),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(net282),
    .B(net384),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _2491_ (.A(net282),
    .B(net384),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _2492_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__o211a_1 _2493_ (.A1(net283),
    .A2(net386),
    .B1(net388),
    .C1(net287),
    .X(_0667_));
 sky130_fd_sc_hd__a21oi_1 _2494_ (.A1(net283),
    .A2(net386),
    .B1(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__o31a_1 _2495_ (.A1(_0654_),
    .A2(_0656_),
    .A3(_0660_),
    .B1(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__or2_1 _2496_ (.A(_0666_),
    .B(net65),
    .X(_0670_));
 sky130_fd_sc_hd__nand2_1 _2497_ (.A(_0666_),
    .B(net65),
    .Y(_0671_));
 sky130_fd_sc_hd__and2_1 _2498_ (.A(_0670_),
    .B(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__or2_1 _2499_ (.A(net456),
    .B(net776),
    .X(_0673_));
 sky130_fd_sc_hd__o211a_1 _2500_ (.A1(net247),
    .A2(_0672_),
    .B1(_0673_),
    .C1(net559),
    .X(_0129_));
 sky130_fd_sc_hd__nand2_1 _2501_ (.A(\scs.acc1[17] ),
    .B(net383),
    .Y(_0674_));
 sky130_fd_sc_hd__inv_2 _2502_ (.A(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _2503_ (.A(\scs.acc1[17] ),
    .B(net383),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _2504_ (.A(_0675_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__a21oi_1 _2505_ (.A1(_0664_),
    .A2(_0670_),
    .B1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__a31o_1 _2506_ (.A1(_0664_),
    .A2(_0670_),
    .A3(_0677_),
    .B1(net249),
    .X(_0679_));
 sky130_fd_sc_hd__nor2_1 _2507_ (.A(net454),
    .B(net382),
    .Y(_0680_));
 sky130_fd_sc_hd__o221a_1 _2508_ (.A1(net455),
    .A2(net383),
    .B1(_0678_),
    .B2(_0679_),
    .C1(net559),
    .X(_0130_));
 sky130_fd_sc_hd__nand2_1 _2509_ (.A(net281),
    .B(net381),
    .Y(_0681_));
 sky130_fd_sc_hd__or2_1 _2510_ (.A(net281),
    .B(net381),
    .X(_0682_));
 sky130_fd_sc_hd__nand2_1 _2511_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a21o_1 _2512_ (.A1(_0664_),
    .A2(_0674_),
    .B1(_0676_),
    .X(_0684_));
 sky130_fd_sc_hd__or3_2 _2513_ (.A(_0666_),
    .B(_0675_),
    .C(_0676_),
    .X(_0685_));
 sky130_fd_sc_hd__o21a_1 _2514_ (.A1(net65),
    .A2(_0685_),
    .B1(_0684_),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_1 _2515_ (.A(_0683_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__or2_1 _2516_ (.A(_0683_),
    .B(_0686_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _2517_ (.A1(_0687_),
    .A2(_0688_),
    .B1(net248),
    .X(_0689_));
 sky130_fd_sc_hd__o211a_1 _2518_ (.A1(net456),
    .A2(net625),
    .B1(net560),
    .C1(_0689_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_1 _2519_ (.A(net279),
    .B(net380),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _2520_ (.A(net279),
    .B(net380),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_1 _2521_ (.A(_0690_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__a21oi_1 _2522_ (.A1(_0681_),
    .A2(_0688_),
    .B1(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__a31o_1 _2523_ (.A1(_0681_),
    .A2(_0688_),
    .A3(_0692_),
    .B1(net247),
    .X(_0694_));
 sky130_fd_sc_hd__o221a_1 _2524_ (.A1(net455),
    .A2(net380),
    .B1(_0693_),
    .B2(_0694_),
    .C1(net559),
    .X(_0132_));
 sky130_fd_sc_hd__nand2_1 _2525_ (.A(\scs.acc1[20] ),
    .B(net378),
    .Y(_0695_));
 sky130_fd_sc_hd__or2_1 _2526_ (.A(\scs.acc1[20] ),
    .B(net378),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _2527_ (.A(_0695_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__or3_1 _2528_ (.A(_0683_),
    .B(_0690_),
    .C(_0691_),
    .X(_0698_));
 sky130_fd_sc_hd__o21ba_1 _2529_ (.A1(_0681_),
    .A2(_0691_),
    .B1_N(_0690_),
    .X(_0699_));
 sky130_fd_sc_hd__o21a_1 _2530_ (.A1(_0684_),
    .A2(_0698_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__o31a_1 _2531_ (.A1(net65),
    .A2(_0685_),
    .A3(_0698_),
    .B1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__xor2_1 _2532_ (.A(_0697_),
    .B(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__or2_1 _2533_ (.A(net460),
    .B(net734),
    .X(_0703_));
 sky130_fd_sc_hd__o211a_1 _2534_ (.A1(net249),
    .A2(_0702_),
    .B1(_0703_),
    .C1(net562),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _2535_ (.A(\scs.acc1[21] ),
    .B(net377),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(\scs.acc1[21] ),
    .B(\scs.acc2[21] ),
    .Y(_0705_));
 sky130_fd_sc_hd__or2_1 _2537_ (.A(_0704_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__o21a_1 _2538_ (.A1(_0697_),
    .A2(_0701_),
    .B1(_0695_),
    .X(_0707_));
 sky130_fd_sc_hd__xnor2_1 _2539_ (.A(_0706_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nor2_1 _2540_ (.A(net457),
    .B(net377),
    .Y(_0709_));
 sky130_fd_sc_hd__a211oi_1 _2541_ (.A1(net457),
    .A2(_0708_),
    .B1(_0709_),
    .C1(net594),
    .Y(_0134_));
 sky130_fd_sc_hd__and2_1 _2542_ (.A(net278),
    .B(net375),
    .X(_0710_));
 sky130_fd_sc_hd__nand2_1 _2543_ (.A(net278),
    .B(net375),
    .Y(_0711_));
 sky130_fd_sc_hd__nor2_1 _2544_ (.A(\scs.acc1[22] ),
    .B(net376),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2_1 _2545_ (.A(_0710_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__or2_1 _2546_ (.A(_0697_),
    .B(_0706_),
    .X(_0714_));
 sky130_fd_sc_hd__o21ba_1 _2547_ (.A1(_0695_),
    .A2(_0705_),
    .B1_N(_0704_),
    .X(_0715_));
 sky130_fd_sc_hd__o21ai_1 _2548_ (.A1(_0701_),
    .A2(_0714_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_1 _2549_ (.A(_0713_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__xnor2_1 _2550_ (.A(_0713_),
    .B(_0716_),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_1 _2551_ (.A(net461),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__o211a_1 _2552_ (.A1(net460),
    .A2(net376),
    .B1(net562),
    .C1(_0719_),
    .X(_0135_));
 sky130_fd_sc_hd__xor2_1 _2553_ (.A(net276),
    .B(net373),
    .X(_0720_));
 sky130_fd_sc_hd__a21oi_1 _2554_ (.A1(_0711_),
    .A2(_0717_),
    .B1(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__a31o_1 _2555_ (.A1(_0711_),
    .A2(_0717_),
    .A3(_0720_),
    .B1(net249),
    .X(_0722_));
 sky130_fd_sc_hd__o221a_1 _2556_ (.A1(net460),
    .A2(net374),
    .B1(_0721_),
    .B2(_0722_),
    .C1(net562),
    .X(_0136_));
 sky130_fd_sc_hd__o21a_1 _2557_ (.A1(_0700_),
    .A2(_0714_),
    .B1(_0715_),
    .X(_0723_));
 sky130_fd_sc_hd__nor2_1 _2558_ (.A(_0712_),
    .B(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a211o_1 _2559_ (.A1(net276),
    .A2(net374),
    .B1(_0710_),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__o21ai_1 _2560_ (.A1(net276),
    .A2(net374),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__or4b_1 _2561_ (.A(_0710_),
    .B(_0712_),
    .C(_0714_),
    .D_N(_0720_),
    .X(_0727_));
 sky130_fd_sc_hd__o41a_1 _2562_ (.A1(_0669_),
    .A2(_0685_),
    .A3(_0698_),
    .A4(_0727_),
    .B1(_0726_),
    .X(_0728_));
 sky130_fd_sc_hd__nand2_1 _2563_ (.A(net275),
    .B(net371),
    .Y(_0729_));
 sky130_fd_sc_hd__or2_1 _2564_ (.A(net275),
    .B(net372),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(_0729_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__xor2_1 _2566_ (.A(_0728_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__or2_1 _2567_ (.A(net468),
    .B(net372),
    .X(_0733_));
 sky130_fd_sc_hd__o211a_1 _2568_ (.A1(net251),
    .A2(_0732_),
    .B1(_0733_),
    .C1(net570),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_1 _2569_ (.A(net274),
    .B(net369),
    .Y(_0734_));
 sky130_fd_sc_hd__inv_2 _2570_ (.A(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2571_ (.A(net274),
    .B(net370),
    .Y(_0736_));
 sky130_fd_sc_hd__nor2_1 _2572_ (.A(_0735_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__o21a_1 _2573_ (.A1(_0728_),
    .A2(_0731_),
    .B1(_0729_),
    .X(_0738_));
 sky130_fd_sc_hd__and2_1 _2574_ (.A(_0737_),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__o21ai_1 _2575_ (.A1(_0737_),
    .A2(_0738_),
    .B1(net464),
    .Y(_0740_));
 sky130_fd_sc_hd__o221a_1 _2576_ (.A1(net464),
    .A2(net370),
    .B1(_0739_),
    .B2(_0740_),
    .C1(net566),
    .X(_0138_));
 sky130_fd_sc_hd__nand2_1 _2577_ (.A(\scs.acc1[26] ),
    .B(net368),
    .Y(_0741_));
 sky130_fd_sc_hd__or2_1 _2578_ (.A(\scs.acc1[26] ),
    .B(net368),
    .X(_0742_));
 sky130_fd_sc_hd__nand2_1 _2579_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__a21o_1 _2580_ (.A1(_0734_),
    .A2(_0738_),
    .B1(_0736_),
    .X(_0744_));
 sky130_fd_sc_hd__or2_1 _2581_ (.A(_0743_),
    .B(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__xnor2_1 _2582_ (.A(_0743_),
    .B(_0744_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _2583_ (.A(net464),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__o211a_1 _2584_ (.A1(net464),
    .A2(net623),
    .B1(net566),
    .C1(_0747_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(\scs.acc1[27] ),
    .B(net367),
    .Y(_0748_));
 sky130_fd_sc_hd__inv_2 _2586_ (.A(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nor2_1 _2587_ (.A(\scs.acc1[27] ),
    .B(net367),
    .Y(_0750_));
 sky130_fd_sc_hd__inv_2 _2588_ (.A(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__o2bb2a_1 _2589_ (.A1_N(_0741_),
    .A2_N(_0745_),
    .B1(_0749_),
    .B2(_0750_),
    .X(_0752_));
 sky130_fd_sc_hd__a41o_1 _2590_ (.A1(_0741_),
    .A2(_0745_),
    .A3(_0748_),
    .A4(_0751_),
    .B1(net251),
    .X(_0753_));
 sky130_fd_sc_hd__o221a_1 _2591_ (.A1(net468),
    .A2(net367),
    .B1(_0752_),
    .B2(_0753_),
    .C1(net570),
    .X(_0140_));
 sky130_fd_sc_hd__or3_1 _2592_ (.A(_0743_),
    .B(_0749_),
    .C(_0750_),
    .X(_0754_));
 sky130_fd_sc_hd__or3_1 _2593_ (.A(_0731_),
    .B(_0735_),
    .C(_0736_),
    .X(_0755_));
 sky130_fd_sc_hd__or3_4 _2594_ (.A(_0728_),
    .B(_0754_),
    .C(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__a211o_1 _2595_ (.A1(_0729_),
    .A2(_0734_),
    .B1(_0736_),
    .C1(_0754_),
    .X(_0757_));
 sky130_fd_sc_hd__or2_1 _2596_ (.A(_0741_),
    .B(_0750_),
    .X(_0758_));
 sky130_fd_sc_hd__and4_1 _2597_ (.A(_0748_),
    .B(_0756_),
    .C(_0757_),
    .D(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _2598_ (.A(net273),
    .B(net365),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _2599_ (.A(net273),
    .B(\scs.acc2[28] ),
    .Y(_0761_));
 sky130_fd_sc_hd__and2b_1 _2600_ (.A_N(_0760_),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__nand2_1 _2601_ (.A(_0759_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21a_1 _2602_ (.A1(_0759_),
    .A2(_0762_),
    .B1(net465),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_1 _2603_ (.A(net465),
    .B(net365),
    .Y(_0765_));
 sky130_fd_sc_hd__a211oi_1 _2604_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0765_),
    .C1(net599),
    .Y(_0141_));
 sky130_fd_sc_hd__a41o_1 _2605_ (.A1(_0748_),
    .A2(_0756_),
    .A3(_0757_),
    .A4(_0758_),
    .B1(_0760_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _2606_ (.A(\scs.acc1[29] ),
    .B(net364),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _2607_ (.A(\scs.acc1[29] ),
    .B(\scs.acc2[29] ),
    .Y(_0768_));
 sky130_fd_sc_hd__and2b_1 _2608_ (.A_N(_0767_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__and3_1 _2609_ (.A(_0761_),
    .B(_0766_),
    .C(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__a21oi_1 _2610_ (.A1(_0761_),
    .A2(_0766_),
    .B1(_0769_),
    .Y(_0771_));
 sky130_fd_sc_hd__or2_1 _2611_ (.A(net465),
    .B(net364),
    .X(_0772_));
 sky130_fd_sc_hd__o311a_1 _2612_ (.A1(net251),
    .A2(_0770_),
    .A3(_0771_),
    .B1(_0772_),
    .C1(net568),
    .X(_0142_));
 sky130_fd_sc_hd__and2_1 _2613_ (.A(net250),
    .B(net363),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_1 _2614_ (.A(net272),
    .B(net363),
    .Y(_0774_));
 sky130_fd_sc_hd__or2_1 _2615_ (.A(net272),
    .B(\scs.acc2[30] ),
    .X(_0775_));
 sky130_fd_sc_hd__and2_1 _2616_ (.A(_0774_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a21o_1 _2617_ (.A1(_0761_),
    .A2(_0766_),
    .B1(_0767_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _2618_ (.A(_0768_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21bo_1 _2619_ (.A1(_0768_),
    .A2(_0777_),
    .B1_N(_0776_),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _2620_ (.A(net468),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o21a_1 _2621_ (.A1(_0776_),
    .A2(_0778_),
    .B1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__o21a_1 _2622_ (.A1(_0773_),
    .A2(_0781_),
    .B1(net568),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _2623_ (.A1(_0774_),
    .A2(_0779_),
    .B1(net468),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _2624_ (.A(net469),
    .B(net655),
    .Y(_0783_));
 sky130_fd_sc_hd__a21oi_1 _2625_ (.A1(_0774_),
    .A2(_0779_),
    .B1(_1475_),
    .Y(_0784_));
 sky130_fd_sc_hd__and3_1 _2626_ (.A(_1475_),
    .B(_0774_),
    .C(_0779_),
    .X(_0785_));
 sky130_fd_sc_hd__o211a_1 _2627_ (.A1(_0784_),
    .A2(_0785_),
    .B1(_0782_),
    .C1(_0783_),
    .X(_0786_));
 sky130_fd_sc_hd__a211o_1 _2628_ (.A1(_0782_),
    .A2(_0783_),
    .B1(_0784_),
    .C1(_0785_),
    .X(_0787_));
 sky130_fd_sc_hd__nor3b_1 _2629_ (.A(net605),
    .B(_0786_),
    .C_N(_0787_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_1 _2630_ (.A1(net435),
    .A2(net412),
    .B1(net361),
    .Y(_0788_));
 sky130_fd_sc_hd__a31o_1 _2631_ (.A1(net435),
    .A2(net876),
    .A3(net412),
    .B1(net582),
    .X(_0789_));
 sky130_fd_sc_hd__nor2_1 _2632_ (.A(_0788_),
    .B(_0789_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand2_1 _2633_ (.A(net359),
    .B(net411),
    .Y(_0790_));
 sky130_fd_sc_hd__or2_1 _2634_ (.A(net360),
    .B(net411),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _2635_ (.A(net362),
    .B(net412),
    .X(_0792_));
 sky130_fd_sc_hd__and3_1 _2636_ (.A(_0790_),
    .B(_0791_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a21oi_1 _2637_ (.A1(_0790_),
    .A2(_0791_),
    .B1(_0792_),
    .Y(_0794_));
 sky130_fd_sc_hd__o21ai_1 _2638_ (.A1(_0793_),
    .A2(_0794_),
    .B1(net434),
    .Y(_0795_));
 sky130_fd_sc_hd__o211a_1 _2639_ (.A1(net434),
    .A2(net360),
    .B1(net515),
    .C1(_0795_),
    .X(_0146_));
 sky130_fd_sc_hd__nor2_1 _2640_ (.A(net358),
    .B(net409),
    .Y(_0796_));
 sky130_fd_sc_hd__and2_1 _2641_ (.A(net812),
    .B(net409),
    .X(_0797_));
 sky130_fd_sc_hd__or2_1 _2642_ (.A(_0796_),
    .B(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a21boi_1 _2643_ (.A1(_0791_),
    .A2(_0792_),
    .B1_N(_0790_),
    .Y(_0799_));
 sky130_fd_sc_hd__a21o_1 _2644_ (.A1(net434),
    .A2(_0799_),
    .B1(_0572_),
    .X(_0800_));
 sky130_fd_sc_hd__a21oi_1 _2645_ (.A1(_0798_),
    .A2(_0800_),
    .B1(net582),
    .Y(_0801_));
 sky130_fd_sc_hd__o31a_1 _2646_ (.A1(_0796_),
    .A2(_0797_),
    .A3(_0800_),
    .B1(_0801_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _2647_ (.A(net357),
    .B(net407),
    .Y(_0802_));
 sky130_fd_sc_hd__and2_1 _2648_ (.A(net814),
    .B(net407),
    .X(_0803_));
 sky130_fd_sc_hd__or2_1 _2649_ (.A(_0802_),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__o21ba_1 _2650_ (.A1(_0796_),
    .A2(_0799_),
    .B1_N(_0797_),
    .X(_0805_));
 sky130_fd_sc_hd__a21o_1 _2651_ (.A1(net438),
    .A2(_0805_),
    .B1(_0579_),
    .X(_0806_));
 sky130_fd_sc_hd__a21oi_1 _2652_ (.A1(_0804_),
    .A2(_0806_),
    .B1(net578),
    .Y(_0807_));
 sky130_fd_sc_hd__o31a_1 _2653_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0806_),
    .B1(_0807_),
    .X(_0148_));
 sky130_fd_sc_hd__o21bai_2 _2654_ (.A1(_0802_),
    .A2(_0805_),
    .B1_N(_0803_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _2655_ (.A(net356),
    .B(net405),
    .Y(_0809_));
 sky130_fd_sc_hd__or2_1 _2656_ (.A(net356),
    .B(net405),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _2657_ (.A(_0809_),
    .B(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _2658_ (.A(_0808_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__or2_1 _2659_ (.A(_0808_),
    .B(_0811_),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _2660_ (.A(_0812_),
    .B(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__or2_1 _2661_ (.A(net430),
    .B(net356),
    .X(_0815_));
 sky130_fd_sc_hd__o211a_1 _2662_ (.A1(net237),
    .A2(_0814_),
    .B1(_0815_),
    .C1(net510),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _2663_ (.A(net354),
    .B(net403),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _2664_ (.A(net354),
    .B(net403),
    .X(_0817_));
 sky130_fd_sc_hd__nand2_1 _2665_ (.A(net353),
    .B(net403),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _2666_ (.A(_0816_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _2667_ (.A(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a31o_1 _2668_ (.A1(net430),
    .A2(_0809_),
    .A3(_0812_),
    .B1(_0593_),
    .X(_0821_));
 sky130_fd_sc_hd__a21oi_1 _2669_ (.A1(_0819_),
    .A2(_0821_),
    .B1(net579),
    .Y(_0822_));
 sky130_fd_sc_hd__o21a_1 _2670_ (.A1(_0819_),
    .A2(_0821_),
    .B1(_0822_),
    .X(_0150_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(net352),
    .B(net401),
    .Y(_0823_));
 sky130_fd_sc_hd__or2_1 _2672_ (.A(net352),
    .B(net401),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _2673_ (.A(_0823_),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _2674_ (.A(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a31o_1 _2675_ (.A1(net356),
    .A2(net405),
    .A3(_0816_),
    .B1(_0817_),
    .X(_0827_));
 sky130_fd_sc_hd__a31o_1 _2676_ (.A1(_0808_),
    .A2(_0811_),
    .A3(_0820_),
    .B1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__nand2_1 _2677_ (.A(_0826_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__xnor2_1 _2678_ (.A(_0825_),
    .B(_0828_),
    .Y(_0830_));
 sky130_fd_sc_hd__or2_1 _2679_ (.A(net430),
    .B(net352),
    .X(_0831_));
 sky130_fd_sc_hd__o211a_1 _2680_ (.A1(net236),
    .A2(_0830_),
    .B1(_0831_),
    .C1(net516),
    .X(_0151_));
 sky130_fd_sc_hd__or2_1 _2681_ (.A(net350),
    .B(net399),
    .X(_0832_));
 sky130_fd_sc_hd__and2_1 _2682_ (.A(net350),
    .B(net399),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _2683_ (.A(net350),
    .B(net399),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _2684_ (.A(_0832_),
    .B(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_2 _2685_ (.A(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__a31o_1 _2686_ (.A1(net432),
    .A2(_0823_),
    .A3(_0829_),
    .B1(_0609_),
    .X(_0837_));
 sky130_fd_sc_hd__a21oi_1 _2687_ (.A1(_0835_),
    .A2(_0837_),
    .B1(net579),
    .Y(_0838_));
 sky130_fd_sc_hd__o21a_1 _2688_ (.A1(_0835_),
    .A2(_0837_),
    .B1(_0838_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _2689_ (.A(net347),
    .B(net397),
    .Y(_0839_));
 sky130_fd_sc_hd__or2_1 _2690_ (.A(net348),
    .B(net397),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_1 _2691_ (.A(_0839_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _2692_ (.A(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a31o_1 _2693_ (.A1(net352),
    .A2(net401),
    .A3(_0832_),
    .B1(_0833_),
    .X(_0843_));
 sky130_fd_sc_hd__a31o_1 _2694_ (.A1(_0826_),
    .A2(_0828_),
    .A3(_0836_),
    .B1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _2695_ (.A(_0842_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__xnor2_1 _2696_ (.A(_0841_),
    .B(_0844_),
    .Y(_0846_));
 sky130_fd_sc_hd__or2_1 _2697_ (.A(net441),
    .B(net348),
    .X(_0847_));
 sky130_fd_sc_hd__o211a_1 _2698_ (.A1(net243),
    .A2(_0846_),
    .B1(_0847_),
    .C1(net516),
    .X(_0153_));
 sky130_fd_sc_hd__or2_1 _2699_ (.A(net346),
    .B(net395),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _2700_ (.A(net346),
    .B(net395),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_2 _2701_ (.A(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _2702_ (.A(_0848_),
    .B(_0849_),
    .Y(_0851_));
 sky130_fd_sc_hd__inv_2 _2703_ (.A(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__a31o_1 _2704_ (.A1(net441),
    .A2(_0839_),
    .A3(_0845_),
    .B1(_0623_),
    .X(_0853_));
 sky130_fd_sc_hd__a21oi_1 _2705_ (.A1(_0851_),
    .A2(_0853_),
    .B1(net586),
    .Y(_0854_));
 sky130_fd_sc_hd__o21a_1 _2706_ (.A1(_0851_),
    .A2(_0853_),
    .B1(_0854_),
    .X(_0154_));
 sky130_fd_sc_hd__nand2_1 _2707_ (.A(net343),
    .B(net394),
    .Y(_0855_));
 sky130_fd_sc_hd__or2_1 _2708_ (.A(net344),
    .B(net394),
    .X(_0856_));
 sky130_fd_sc_hd__a31o_1 _2709_ (.A1(net348),
    .A2(net397),
    .A3(_0848_),
    .B1(_0850_),
    .X(_0857_));
 sky130_fd_sc_hd__a31o_1 _2710_ (.A1(_0842_),
    .A2(_0844_),
    .A3(_0852_),
    .B1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__a21o_1 _2711_ (.A1(_0855_),
    .A2(_0856_),
    .B1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__nand3_1 _2712_ (.A(_0855_),
    .B(_0856_),
    .C(_0858_),
    .Y(_0860_));
 sky130_fd_sc_hd__and3_1 _2713_ (.A(net441),
    .B(_0859_),
    .C(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__a21oi_1 _2714_ (.A1(net243),
    .A2(net344),
    .B1(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(net588),
    .B(_0862_),
    .Y(_0155_));
 sky130_fd_sc_hd__and2_1 _2716_ (.A(net341),
    .B(net393),
    .X(_0863_));
 sky130_fd_sc_hd__or2_1 _2717_ (.A(net342),
    .B(net393),
    .X(_0864_));
 sky130_fd_sc_hd__nand2b_1 _2718_ (.A_N(_0863_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__a21bo_1 _2719_ (.A1(_0856_),
    .A2(_0858_),
    .B1_N(_0855_),
    .X(_0866_));
 sky130_fd_sc_hd__xnor2_1 _2720_ (.A(_0865_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(net342),
    .A1(_0867_),
    .S(net443),
    .X(_0868_));
 sky130_fd_sc_hd__and2_1 _2722_ (.A(net517),
    .B(_0868_),
    .X(_0156_));
 sky130_fd_sc_hd__a21oi_2 _2723_ (.A1(_0864_),
    .A2(_0866_),
    .B1(_0863_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _2724_ (.A(net340),
    .B(net391),
    .Y(_0870_));
 sky130_fd_sc_hd__or2_1 _2725_ (.A(net340),
    .B(net391),
    .X(_0871_));
 sky130_fd_sc_hd__nand2_1 _2726_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__or2_1 _2727_ (.A(_0869_),
    .B(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__xor2_1 _2728_ (.A(_0869_),
    .B(_0872_),
    .X(_0874_));
 sky130_fd_sc_hd__or2_1 _2729_ (.A(net443),
    .B(net340),
    .X(_0875_));
 sky130_fd_sc_hd__o211a_1 _2730_ (.A1(net244),
    .A2(_0874_),
    .B1(_0875_),
    .C1(net518),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _2731_ (.A(net337),
    .B(net389),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_1 _2732_ (.A(net338),
    .B(net389),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_1 _2733_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__a31o_1 _2734_ (.A1(net443),
    .A2(_0870_),
    .A3(_0873_),
    .B1(_0651_),
    .X(_0879_));
 sky130_fd_sc_hd__a21oi_1 _2735_ (.A1(_0878_),
    .A2(_0879_),
    .B1(net588),
    .Y(_0880_));
 sky130_fd_sc_hd__o21a_1 _2736_ (.A1(_0878_),
    .A2(_0879_),
    .B1(_0880_),
    .X(_0158_));
 sky130_fd_sc_hd__nand2_1 _2737_ (.A(net336),
    .B(net387),
    .Y(_0881_));
 sky130_fd_sc_hd__or2_1 _2738_ (.A(net336),
    .B(net387),
    .X(_0882_));
 sky130_fd_sc_hd__nand2_1 _2739_ (.A(_0881_),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__and3_1 _2740_ (.A(net340),
    .B(net391),
    .C(_0876_),
    .X(_0884_));
 sky130_fd_sc_hd__a21oi_1 _2741_ (.A1(net338),
    .A2(net389),
    .B1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__o31a_1 _2742_ (.A1(_0869_),
    .A2(_0872_),
    .A3(_0878_),
    .B1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or2_1 _2743_ (.A(_0883_),
    .B(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__xor2_1 _2744_ (.A(_0883_),
    .B(_0886_),
    .X(_0888_));
 sky130_fd_sc_hd__or2_1 _2745_ (.A(net444),
    .B(net336),
    .X(_0889_));
 sky130_fd_sc_hd__o211a_1 _2746_ (.A1(net244),
    .A2(_0888_),
    .B1(_0889_),
    .C1(net558),
    .X(_0159_));
 sky130_fd_sc_hd__xnor2_1 _2747_ (.A(net333),
    .B(net385),
    .Y(_0890_));
 sky130_fd_sc_hd__a31o_1 _2748_ (.A1(net444),
    .A2(_0881_),
    .A3(_0887_),
    .B1(_0663_),
    .X(_0891_));
 sky130_fd_sc_hd__a21oi_1 _2749_ (.A1(_0890_),
    .A2(_0891_),
    .B1(net594),
    .Y(_0892_));
 sky130_fd_sc_hd__o21a_1 _2750_ (.A1(_0890_),
    .A2(_0891_),
    .B1(_0892_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _2751_ (.A(net331),
    .B(net384),
    .Y(_0893_));
 sky130_fd_sc_hd__or2_1 _2752_ (.A(net332),
    .B(net384),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _2753_ (.A(_0893_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__o211a_1 _2754_ (.A1(net334),
    .A2(net385),
    .B1(net387),
    .C1(net336),
    .X(_0896_));
 sky130_fd_sc_hd__a21oi_1 _2755_ (.A1(net334),
    .A2(net385),
    .B1(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__o31a_1 _2756_ (.A1(_0883_),
    .A2(_0886_),
    .A3(_0890_),
    .B1(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__or2_1 _2757_ (.A(_0895_),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _2758_ (.A(_0895_),
    .B(_0898_),
    .Y(_0900_));
 sky130_fd_sc_hd__and2_1 _2759_ (.A(_0899_),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__or2_1 _2760_ (.A(net454),
    .B(net332),
    .X(_0902_));
 sky130_fd_sc_hd__o211a_1 _2761_ (.A1(net247),
    .A2(_0901_),
    .B1(_0902_),
    .C1(net558),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _2762_ (.A(net330),
    .B(net382),
    .Y(_0903_));
 sky130_fd_sc_hd__nor2_1 _2763_ (.A(net330),
    .B(net382),
    .Y(_0904_));
 sky130_fd_sc_hd__or2_1 _2764_ (.A(net330),
    .B(net382),
    .X(_0905_));
 sky130_fd_sc_hd__nand2_1 _2765_ (.A(_0903_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__a31o_1 _2766_ (.A1(net454),
    .A2(_0893_),
    .A3(_0899_),
    .B1(_0680_),
    .X(_0907_));
 sky130_fd_sc_hd__a21oi_1 _2767_ (.A1(_0906_),
    .A2(_0907_),
    .B1(net594),
    .Y(_0908_));
 sky130_fd_sc_hd__o21a_1 _2768_ (.A1(_0906_),
    .A2(_0907_),
    .B1(_0908_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _2769_ (.A(net247),
    .B(net327),
    .Y(_0909_));
 sky130_fd_sc_hd__and2_1 _2770_ (.A(net328),
    .B(net381),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_1 _2771_ (.A(net328),
    .B(net381),
    .Y(_0911_));
 sky130_fd_sc_hd__or2_1 _2772_ (.A(_0910_),
    .B(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__a31o_1 _2773_ (.A1(_0893_),
    .A2(_0899_),
    .A3(_0903_),
    .B1(_0904_),
    .X(_0913_));
 sky130_fd_sc_hd__o21ai_1 _2774_ (.A1(_0912_),
    .A2(_0913_),
    .B1(net454),
    .Y(_0914_));
 sky130_fd_sc_hd__a21o_1 _2775_ (.A1(_0912_),
    .A2(_0913_),
    .B1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a21oi_1 _2776_ (.A1(_0909_),
    .A2(_0915_),
    .B1(net595),
    .Y(_0163_));
 sky130_fd_sc_hd__and2_1 _2777_ (.A(net325),
    .B(net379),
    .X(_0916_));
 sky130_fd_sc_hd__nor2_1 _2778_ (.A(net326),
    .B(net379),
    .Y(_0917_));
 sky130_fd_sc_hd__or2_1 _2779_ (.A(net326),
    .B(net379),
    .X(_0918_));
 sky130_fd_sc_hd__or2_1 _2780_ (.A(_0916_),
    .B(_0917_),
    .X(_0919_));
 sky130_fd_sc_hd__o22ai_1 _2781_ (.A1(net455),
    .A2(net379),
    .B1(_0910_),
    .B2(_0914_),
    .Y(_0920_));
 sky130_fd_sc_hd__xnor2_1 _2782_ (.A(_0919_),
    .B(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2_1 _2783_ (.A(net595),
    .B(_0921_),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_1 _2784_ (.A(net323),
    .B(net378),
    .Y(_0922_));
 sky130_fd_sc_hd__or2_1 _2785_ (.A(net324),
    .B(net378),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _2786_ (.A(_0922_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__or3_1 _2787_ (.A(_0912_),
    .B(_0916_),
    .C(_0917_),
    .X(_0925_));
 sky130_fd_sc_hd__or3_1 _2788_ (.A(_0895_),
    .B(_0906_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__a211oi_1 _2789_ (.A1(_0893_),
    .A2(_0903_),
    .B1(_0904_),
    .C1(_0925_),
    .Y(_0927_));
 sky130_fd_sc_hd__a211o_1 _2790_ (.A1(_0910_),
    .A2(_0918_),
    .B1(_0927_),
    .C1(_0916_),
    .X(_0928_));
 sky130_fd_sc_hd__o21ba_1 _2791_ (.A1(_0898_),
    .A2(_0926_),
    .B1_N(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__xor2_1 _2792_ (.A(_0924_),
    .B(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__or2_1 _2793_ (.A(net458),
    .B(net324),
    .X(_0931_));
 sky130_fd_sc_hd__o211a_1 _2794_ (.A1(net248),
    .A2(_0930_),
    .B1(_0931_),
    .C1(net561),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_1 _2795_ (.A(net322),
    .B(net377),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _2796_ (.A(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_1 _2797_ (.A(net322),
    .B(net377),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_1 _2798_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__o21a_1 _2799_ (.A1(_0924_),
    .A2(_0929_),
    .B1(_0922_),
    .X(_0936_));
 sky130_fd_sc_hd__a21oi_1 _2800_ (.A1(net457),
    .A2(_0936_),
    .B1(_0709_),
    .Y(_0937_));
 sky130_fd_sc_hd__xnor2_1 _2801_ (.A(_0935_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_1 _2802_ (.A(net595),
    .B(_0938_),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _2803_ (.A(net248),
    .B(net319),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _2804_ (.A(net320),
    .B(net375),
    .Y(_0940_));
 sky130_fd_sc_hd__or2_1 _2805_ (.A(net320),
    .B(net375),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _2806_ (.A(_0940_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__a21o_1 _2807_ (.A1(_0932_),
    .A2(_0936_),
    .B1(_0934_),
    .X(_0943_));
 sky130_fd_sc_hd__o21a_1 _2808_ (.A1(_0942_),
    .A2(_0943_),
    .B1(net457),
    .X(_0944_));
 sky130_fd_sc_hd__a21bo_1 _2809_ (.A1(_0942_),
    .A2(_0943_),
    .B1_N(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__a21oi_1 _2810_ (.A1(_0939_),
    .A2(_0945_),
    .B1(net600),
    .Y(_0167_));
 sky130_fd_sc_hd__or2_1 _2811_ (.A(net318),
    .B(net373),
    .X(_0946_));
 sky130_fd_sc_hd__nand2_1 _2812_ (.A(\scs.acc3[23] ),
    .B(net373),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _2813_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a2bb2o_1 _2814_ (.A1_N(net458),
    .A2_N(net373),
    .B1(_0940_),
    .B2(_0944_),
    .X(_0949_));
 sky130_fd_sc_hd__a21oi_1 _2815_ (.A1(_0948_),
    .A2(_0949_),
    .B1(net600),
    .Y(_0950_));
 sky130_fd_sc_hd__o21a_1 _2816_ (.A1(_0948_),
    .A2(_0949_),
    .B1(_0950_),
    .X(_0168_));
 sky130_fd_sc_hd__nand2_1 _2817_ (.A(net316),
    .B(net371),
    .Y(_0951_));
 sky130_fd_sc_hd__or2_1 _2818_ (.A(net317),
    .B(net371),
    .X(_0952_));
 sky130_fd_sc_hd__nand2_1 _2819_ (.A(_0951_),
    .B(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__or4_1 _2820_ (.A(_0924_),
    .B(_0933_),
    .C(_0934_),
    .D(_0942_),
    .X(_0954_));
 sky130_fd_sc_hd__or2_1 _2821_ (.A(_0948_),
    .B(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o21a_1 _2822_ (.A1(_0922_),
    .A2(_0934_),
    .B1(_0932_),
    .X(_0956_));
 sky130_fd_sc_hd__a21bo_1 _2823_ (.A1(_0940_),
    .A2(_0947_),
    .B1_N(_0946_),
    .X(_0957_));
 sky130_fd_sc_hd__nand2b_1 _2824_ (.A_N(_0955_),
    .B(_0928_),
    .Y(_0958_));
 sky130_fd_sc_hd__o311a_1 _2825_ (.A1(_0942_),
    .A2(_0948_),
    .A3(_0956_),
    .B1(_0957_),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__o31a_1 _2826_ (.A1(_0898_),
    .A2(_0926_),
    .A3(_0955_),
    .B1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__or2_1 _2827_ (.A(_0953_),
    .B(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__nand2_1 _2828_ (.A(_0953_),
    .B(_0960_),
    .Y(_0962_));
 sky130_fd_sc_hd__and2_1 _2829_ (.A(_0961_),
    .B(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2830_ (.A(net463),
    .B(net317),
    .X(_0964_));
 sky130_fd_sc_hd__o211a_1 _2831_ (.A1(net250),
    .A2(_0963_),
    .B1(_0964_),
    .C1(net564),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _2832_ (.A(net315),
    .B(net369),
    .X(_0965_));
 sky130_fd_sc_hd__nor2_1 _2833_ (.A(\scs.acc3[25] ),
    .B(net369),
    .Y(_0966_));
 sky130_fd_sc_hd__or2_1 _2834_ (.A(_0965_),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(_0951_),
    .B(_0961_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(net369),
    .A1(_0968_),
    .S(net463),
    .X(_0969_));
 sky130_fd_sc_hd__xor2_1 _2837_ (.A(_0967_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_1 _2838_ (.A(net600),
    .B(_0970_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_1 _2839_ (.A(net313),
    .B(net368),
    .Y(_0971_));
 sky130_fd_sc_hd__or2_1 _2840_ (.A(net314),
    .B(net368),
    .X(_0972_));
 sky130_fd_sc_hd__nand2_1 _2841_ (.A(_0971_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__o21bai_1 _2842_ (.A1(_0965_),
    .A2(_0968_),
    .B1_N(_0966_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _2843_ (.A(_0973_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__o21a_1 _2844_ (.A1(_0973_),
    .A2(_0974_),
    .B1(net463),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _2845_ (.A1(net250),
    .A2(net314),
    .B1(_0975_),
    .B2(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__and2_1 _2846_ (.A(net565),
    .B(_0977_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _2847_ (.A(net312),
    .B(net366),
    .Y(_0978_));
 sky130_fd_sc_hd__nor2_1 _2848_ (.A(net312),
    .B(net366),
    .Y(_0979_));
 sky130_fd_sc_hd__or2_1 _2849_ (.A(net311),
    .B(net366),
    .X(_0980_));
 sky130_fd_sc_hd__nand2_1 _2850_ (.A(_0978_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__a2bb2o_1 _2851_ (.A1_N(net463),
    .A2_N(net366),
    .B1(_0971_),
    .B2(_0976_),
    .X(_0982_));
 sky130_fd_sc_hd__a21oi_1 _2852_ (.A1(_0981_),
    .A2(_0982_),
    .B1(net599),
    .Y(_0983_));
 sky130_fd_sc_hd__o21a_1 _2853_ (.A1(_0981_),
    .A2(_0982_),
    .B1(_0983_),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_1 _2854_ (.A(net310),
    .B(net365),
    .Y(_0984_));
 sky130_fd_sc_hd__and2_1 _2855_ (.A(net850),
    .B(net365),
    .X(_0985_));
 sky130_fd_sc_hd__or2_1 _2856_ (.A(_0984_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__or3_1 _2857_ (.A(_0967_),
    .B(_0973_),
    .C(_0981_),
    .X(_0987_));
 sky130_fd_sc_hd__a21oi_1 _2858_ (.A1(net317),
    .A2(net371),
    .B1(_0965_),
    .Y(_0988_));
 sky130_fd_sc_hd__or4_1 _2859_ (.A(_0966_),
    .B(_0973_),
    .C(_0981_),
    .D(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__o211a_1 _2860_ (.A1(_0971_),
    .A2(_0979_),
    .B1(_0989_),
    .C1(_0978_),
    .X(_0990_));
 sky130_fd_sc_hd__o21a_1 _2861_ (.A1(_0961_),
    .A2(_0987_),
    .B1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__a21o_1 _2862_ (.A1(net466),
    .A2(_0991_),
    .B1(_0765_),
    .X(_0992_));
 sky130_fd_sc_hd__a21oi_1 _2863_ (.A1(_0986_),
    .A2(_0992_),
    .B1(net599),
    .Y(_0993_));
 sky130_fd_sc_hd__o31a_1 _2864_ (.A1(_0984_),
    .A2(_0985_),
    .A3(_0992_),
    .B1(_0993_),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_1 _2865_ (.A(net309),
    .B(net364),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _2866_ (.A(net804),
    .B(net364),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2b_1 _2867_ (.A_N(_0994_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__o21ba_1 _2868_ (.A1(_0984_),
    .A2(_0991_),
    .B1_N(_0985_),
    .X(_0997_));
 sky130_fd_sc_hd__a21bo_1 _2869_ (.A1(net465),
    .A2(_0997_),
    .B1_N(_0772_),
    .X(_0998_));
 sky130_fd_sc_hd__a21oi_1 _2870_ (.A1(_0996_),
    .A2(_0998_),
    .B1(net599),
    .Y(_0999_));
 sky130_fd_sc_hd__o21a_1 _2871_ (.A1(_0996_),
    .A2(_0998_),
    .B1(_0999_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _2872_ (.A(net695),
    .B(net363),
    .Y(_1000_));
 sky130_fd_sc_hd__or2_1 _2873_ (.A(net695),
    .B(net363),
    .X(_1001_));
 sky130_fd_sc_hd__nand2_1 _2874_ (.A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__o21a_1 _2875_ (.A1(_0994_),
    .A2(_0997_),
    .B1(_0995_),
    .X(_1003_));
 sky130_fd_sc_hd__xnor2_1 _2876_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _2877_ (.A(net466),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__o211a_1 _2878_ (.A1(net466),
    .A2(net792),
    .B1(net568),
    .C1(_1005_),
    .X(_0175_));
 sky130_fd_sc_hd__o21a_1 _2879_ (.A1(_1002_),
    .A2(_1003_),
    .B1(_1000_),
    .X(_1006_));
 sky130_fd_sc_hd__xor2_1 _2880_ (.A(\scs.acc3[31] ),
    .B(\scs.acc2[31] ),
    .X(_1007_));
 sky130_fd_sc_hd__xnor2_1 _2881_ (.A(_1006_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__or2_1 _2882_ (.A(net467),
    .B(\scs.acc3[31] ),
    .X(_1009_));
 sky130_fd_sc_hd__o211a_1 _2883_ (.A1(net250),
    .A2(_1008_),
    .B1(_1009_),
    .C1(net568),
    .X(_0176_));
 sky130_fd_sc_hd__xor2_2 _2884_ (.A(\pr.genblk1[1].pd.ff_reg_1 ),
    .B(\pr.genblk1[1].pd.ff_reg_0 ),
    .X(_1010_));
 sky130_fd_sc_hd__xor2_2 _2885_ (.A(\pr.genblk1[0].pd.ff_reg_1 ),
    .B(\pr.genblk1[0].pd.ff_reg_0 ),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_1 _2886_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__xnor2_2 _2887_ (.A(_1010_),
    .B(_1011_),
    .Y(_1013_));
 sky130_fd_sc_hd__xnor2_2 _2888_ (.A(\pr.genblk1[10].pd.ff_reg_1 ),
    .B(\pr.genblk1[10].pd.ff_reg_0 ),
    .Y(_1014_));
 sky130_fd_sc_hd__and2b_1 _2889_ (.A_N(_1013_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__xor2_2 _2890_ (.A(_1013_),
    .B(_1014_),
    .X(_1016_));
 sky130_fd_sc_hd__xor2_4 _2891_ (.A(\pr.genblk1[8].pd.ff_reg_1 ),
    .B(\pr.genblk1[8].pd.ff_reg_0 ),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_1 _2892_ (.A(_1016_),
    .B(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__xnor2_2 _2893_ (.A(_1016_),
    .B(_1017_),
    .Y(_1019_));
 sky130_fd_sc_hd__xnor2_1 _2894_ (.A(\pr.genblk1[3].pd.ff_reg_1 ),
    .B(\pr.genblk1[3].pd.ff_reg_0 ),
    .Y(_1020_));
 sky130_fd_sc_hd__and2b_1 _2895_ (.A_N(_1019_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__xnor2_2 _2896_ (.A(_1019_),
    .B(_1020_),
    .Y(_1022_));
 sky130_fd_sc_hd__xor2_1 _2897_ (.A(\pr.genblk1[6].pd.ff_reg_1 ),
    .B(\pr.genblk1[6].pd.ff_reg_0 ),
    .X(_1023_));
 sky130_fd_sc_hd__or2_1 _2898_ (.A(\pr.genblk1[4].pd.ff_reg_1 ),
    .B(\pr.genblk1[4].pd.ff_reg_0 ),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _2899_ (.A(\pr.genblk1[4].pd.ff_reg_1 ),
    .B(\pr.genblk1[4].pd.ff_reg_0 ),
    .Y(_1025_));
 sky130_fd_sc_hd__a21o_1 _2900_ (.A1(_1024_),
    .A2(_1025_),
    .B1(_1023_),
    .X(_1026_));
 sky130_fd_sc_hd__nand3_1 _2901_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _2902_ (.A(_1026_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__xnor2_2 _2903_ (.A(\pr.genblk1[2].pd.ff_reg_1 ),
    .B(\pr.genblk1[2].pd.ff_reg_0 ),
    .Y(_1029_));
 sky130_fd_sc_hd__xnor2_2 _2904_ (.A(_1028_),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__xnor2_2 _2905_ (.A(_1022_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__xnor2_2 _2906_ (.A(\pr.genblk1[7].pd.ff_reg_1 ),
    .B(\pr.genblk1[7].pd.ff_reg_0 ),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2b_1 _2907_ (.A_N(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__xnor2_2 _2908_ (.A(_1031_),
    .B(_1032_),
    .Y(_1034_));
 sky130_fd_sc_hd__xnor2_2 _2909_ (.A(\pr.genblk1[5].pd.ff_reg_1 ),
    .B(\pr.genblk1[5].pd.ff_reg_0 ),
    .Y(_1035_));
 sky130_fd_sc_hd__xnor2_2 _2910_ (.A(_1034_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__xnor2_2 _2911_ (.A(\pr.genblk1[9].pd.ff_reg_1 ),
    .B(\pr.genblk1[9].pd.ff_reg_0 ),
    .Y(_1037_));
 sky130_fd_sc_hd__and2b_1 _2912_ (.A_N(_1036_),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__xnor2_2 _2913_ (.A(_1036_),
    .B(_1037_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _2914_ (.A(net830),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__a21o_1 _2915_ (.A1(net450),
    .A2(_1039_),
    .B1(net830),
    .X(_1041_));
 sky130_fd_sc_hd__o211a_1 _2916_ (.A1(net241),
    .A2(_1040_),
    .B1(_1041_),
    .C1(net518),
    .X(_0177_));
 sky130_fd_sc_hd__a21bo_1 _2917_ (.A1(_1027_),
    .A2(_1029_),
    .B1_N(_1026_),
    .X(_1042_));
 sky130_fd_sc_hd__a21o_1 _2918_ (.A1(_1022_),
    .A2(_1030_),
    .B1(_1021_),
    .X(_1043_));
 sky130_fd_sc_hd__nand2_1 _2919_ (.A(_1012_),
    .B(_1018_),
    .Y(_1044_));
 sky130_fd_sc_hd__xor2_1 _2920_ (.A(_1012_),
    .B(_1018_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(_1015_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__o21a_1 _2922_ (.A1(_1015_),
    .A2(_1045_),
    .B1(_1043_),
    .X(_1047_));
 sky130_fd_sc_hd__xor2_2 _2923_ (.A(_1043_),
    .B(_1046_),
    .X(_1048_));
 sky130_fd_sc_hd__and2b_1 _2924_ (.A_N(_1048_),
    .B(_1042_),
    .X(_1049_));
 sky130_fd_sc_hd__xor2_2 _2925_ (.A(_1042_),
    .B(_1048_),
    .X(_1050_));
 sky130_fd_sc_hd__a21boi_2 _2926_ (.A1(_1034_),
    .A2(_1035_),
    .B1_N(_1033_),
    .Y(_1051_));
 sky130_fd_sc_hd__nor2_1 _2927_ (.A(_1050_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__xor2_2 _2928_ (.A(_1050_),
    .B(_1051_),
    .X(_1053_));
 sky130_fd_sc_hd__xor2_2 _2929_ (.A(_1038_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _2930_ (.A(net308),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__xnor2_1 _2931_ (.A(\scs.acc1[1] ),
    .B(_1054_),
    .Y(_1056_));
 sky130_fd_sc_hd__xnor2_1 _2932_ (.A(_1040_),
    .B(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(_1471_),
    .A1(_1057_),
    .S(net450),
    .X(_1058_));
 sky130_fd_sc_hd__nor2_1 _2934_ (.A(net589),
    .B(_1058_),
    .Y(_0178_));
 sky130_fd_sc_hd__a21o_1 _2935_ (.A1(_1038_),
    .A2(_1053_),
    .B1(_1052_),
    .X(_1059_));
 sky130_fd_sc_hd__nor2_1 _2936_ (.A(_1047_),
    .B(_1049_),
    .Y(_1060_));
 sky130_fd_sc_hd__nor2_1 _2937_ (.A(_1044_),
    .B(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__xnor2_2 _2938_ (.A(_1044_),
    .B(_1060_),
    .Y(_1062_));
 sky130_fd_sc_hd__and2b_1 _2939_ (.A_N(_1062_),
    .B(_1059_),
    .X(_1063_));
 sky130_fd_sc_hd__xnor2_1 _2940_ (.A(_1059_),
    .B(_1062_),
    .Y(_1064_));
 sky130_fd_sc_hd__and2_1 _2941_ (.A(net306),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__or2_1 _2942_ (.A(net307),
    .B(_1064_),
    .X(_1066_));
 sky130_fd_sc_hd__nand2b_1 _2943_ (.A_N(_1065_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__o21ai_1 _2944_ (.A1(_1040_),
    .A2(_1056_),
    .B1(_1055_),
    .Y(_1068_));
 sky130_fd_sc_hd__xnor2_1 _2945_ (.A(_1067_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(net307),
    .A1(_1069_),
    .S(net449),
    .X(_1070_));
 sky130_fd_sc_hd__and2_1 _2947_ (.A(net519),
    .B(_1070_),
    .X(_0179_));
 sky130_fd_sc_hd__o21a_1 _2948_ (.A1(_1061_),
    .A2(_1063_),
    .B1(net305),
    .X(_1071_));
 sky130_fd_sc_hd__or3_1 _2949_ (.A(net305),
    .B(_1061_),
    .C(_1063_),
    .X(_1072_));
 sky130_fd_sc_hd__nand2b_1 _2950_ (.A_N(_1071_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__a21o_1 _2951_ (.A1(_1066_),
    .A2(_1068_),
    .B1(_1065_),
    .X(_1074_));
 sky130_fd_sc_hd__xnor2_1 _2952_ (.A(_1073_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(net304),
    .A1(_1075_),
    .S(net450),
    .X(_1076_));
 sky130_fd_sc_hd__and2_1 _2954_ (.A(net518),
    .B(_1076_),
    .X(_0180_));
 sky130_fd_sc_hd__a21o_1 _2955_ (.A1(_1072_),
    .A2(_1074_),
    .B1(_1071_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _2956_ (.A(net449),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__inv_2 _2957_ (.A(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__a21oi_1 _2958_ (.A1(net301),
    .A2(_1079_),
    .B1(net584),
    .Y(_1080_));
 sky130_fd_sc_hd__o21a_1 _2959_ (.A1(net301),
    .A2(_1079_),
    .B1(_1080_),
    .X(_0181_));
 sky130_fd_sc_hd__a21oi_1 _2960_ (.A1(net301),
    .A2(_1079_),
    .B1(net300),
    .Y(_1081_));
 sky130_fd_sc_hd__and3_1 _2961_ (.A(\scs.acc1[5] ),
    .B(net301),
    .C(_1079_),
    .X(_1082_));
 sky130_fd_sc_hd__nor3_1 _2962_ (.A(net584),
    .B(_1081_),
    .C(net867),
    .Y(_0182_));
 sky130_fd_sc_hd__a21oi_1 _2963_ (.A1(net299),
    .A2(_1082_),
    .B1(net584),
    .Y(_1083_));
 sky130_fd_sc_hd__o21a_1 _2964_ (.A1(net299),
    .A2(_1082_),
    .B1(_1083_),
    .X(_0183_));
 sky130_fd_sc_hd__a21oi_1 _2965_ (.A1(net298),
    .A2(_1082_),
    .B1(net712),
    .Y(_1084_));
 sky130_fd_sc_hd__and4_1 _2966_ (.A(\scs.acc1[7] ),
    .B(net299),
    .C(net300),
    .D(net302),
    .X(_1085_));
 sky130_fd_sc_hd__and3_1 _2967_ (.A(net449),
    .B(_1077_),
    .C(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__nor3_1 _2968_ (.A(net584),
    .B(_1084_),
    .C(net63),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _2969_ (.A1(net296),
    .A2(net63),
    .B1(net585),
    .Y(_1087_));
 sky130_fd_sc_hd__o21a_1 _2970_ (.A1(net296),
    .A2(net63),
    .B1(_1087_),
    .X(_0185_));
 sky130_fd_sc_hd__a21oi_1 _2971_ (.A1(net296),
    .A2(net63),
    .B1(net294),
    .Y(_1088_));
 sky130_fd_sc_hd__and3_1 _2972_ (.A(net295),
    .B(net296),
    .C(_1086_),
    .X(_1089_));
 sky130_fd_sc_hd__nor3_1 _2973_ (.A(net585),
    .B(_1088_),
    .C(_1089_),
    .Y(_0186_));
 sky130_fd_sc_hd__or2_1 _2974_ (.A(net803),
    .B(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nand2_1 _2975_ (.A(net293),
    .B(_1089_),
    .Y(_1091_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(net519),
    .B(_1090_),
    .C(_1091_),
    .X(_0187_));
 sky130_fd_sc_hd__and4_1 _2977_ (.A(\scs.acc1[11] ),
    .B(net293),
    .C(net295),
    .D(\scs.acc1[8] ),
    .X(_1092_));
 sky130_fd_sc_hd__and4_1 _2978_ (.A(net449),
    .B(_1077_),
    .C(_1085_),
    .D(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__a211oi_1 _2979_ (.A1(_1470_),
    .A2(_1091_),
    .B1(_1093_),
    .C1(net589),
    .Y(_0188_));
 sky130_fd_sc_hd__and2_1 _2980_ (.A(net291),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _2981_ (.A(net589),
    .B(net61),
    .Y(_1095_));
 sky130_fd_sc_hd__o21a_1 _2982_ (.A1(net292),
    .A2(_1093_),
    .B1(_1095_),
    .X(_0189_));
 sky130_fd_sc_hd__a21oi_1 _2983_ (.A1(net288),
    .A2(net61),
    .B1(net589),
    .Y(_1096_));
 sky130_fd_sc_hd__o21a_1 _2984_ (.A1(net288),
    .A2(net61),
    .B1(_1096_),
    .X(_0190_));
 sky130_fd_sc_hd__a21oi_1 _2985_ (.A1(net289),
    .A2(net62),
    .B1(net285),
    .Y(_1097_));
 sky130_fd_sc_hd__a31o_1 _2986_ (.A1(net286),
    .A2(net288),
    .A3(net62),
    .B1(net590),
    .X(_1098_));
 sky130_fd_sc_hd__nor2_1 _2987_ (.A(_1097_),
    .B(_1098_),
    .Y(_0191_));
 sky130_fd_sc_hd__a31oi_1 _2988_ (.A1(net285),
    .A2(net289),
    .A3(net62),
    .B1(net283),
    .Y(_1099_));
 sky130_fd_sc_hd__and4_1 _2989_ (.A(net284),
    .B(net285),
    .C(net289),
    .D(net61),
    .X(_1100_));
 sky130_fd_sc_hd__nor3_1 _2990_ (.A(net596),
    .B(_1099_),
    .C(net59),
    .Y(_0192_));
 sky130_fd_sc_hd__and2_1 _2991_ (.A(net282),
    .B(net57),
    .X(_1101_));
 sky130_fd_sc_hd__nor2_1 _2992_ (.A(net282),
    .B(net57),
    .Y(_1102_));
 sky130_fd_sc_hd__nor3_1 _2993_ (.A(net596),
    .B(_1101_),
    .C(_1102_),
    .Y(_0193_));
 sky130_fd_sc_hd__and2_1 _2994_ (.A(\scs.acc1[17] ),
    .B(\scs.acc1[16] ),
    .X(_1103_));
 sky130_fd_sc_hd__nand2_1 _2995_ (.A(net57),
    .B(net70),
    .Y(_1104_));
 sky130_fd_sc_hd__o211a_1 _2996_ (.A1(net738),
    .A2(_1101_),
    .B1(_1104_),
    .C1(net562),
    .X(_0194_));
 sky130_fd_sc_hd__a21oi_1 _2997_ (.A1(net57),
    .A2(net69),
    .B1(net280),
    .Y(_1105_));
 sky130_fd_sc_hd__a31o_1 _2998_ (.A1(net280),
    .A2(net58),
    .A3(net69),
    .B1(net596),
    .X(_1106_));
 sky130_fd_sc_hd__nor2_1 _2999_ (.A(_1105_),
    .B(_1106_),
    .Y(_0195_));
 sky130_fd_sc_hd__a31oi_1 _3000_ (.A1(net280),
    .A2(net58),
    .A3(net69),
    .B1(net279),
    .Y(_1107_));
 sky130_fd_sc_hd__and4_1 _3001_ (.A(net279),
    .B(net280),
    .C(net58),
    .D(net70),
    .X(_1108_));
 sky130_fd_sc_hd__nor3_1 _3002_ (.A(net596),
    .B(_1107_),
    .C(_1108_),
    .Y(_0196_));
 sky130_fd_sc_hd__and3_1 _3003_ (.A(\scs.acc1[19] ),
    .B(net281),
    .C(net69),
    .X(_1109_));
 sky130_fd_sc_hd__and3_1 _3004_ (.A(net460),
    .B(\scs.acc1[20] ),
    .C(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__and4_1 _3005_ (.A(net284),
    .B(net285),
    .C(net288),
    .D(net292),
    .X(_1111_));
 sky130_fd_sc_hd__and4_1 _3006_ (.A(_1077_),
    .B(_1085_),
    .C(_1092_),
    .D(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__nand2_1 _3007_ (.A(_1110_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__o211a_1 _3008_ (.A1(net711),
    .A2(_1108_),
    .B1(_1113_),
    .C1(net563),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_1 _3009_ (.A(_1469_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__xnor2_1 _3010_ (.A(_1469_),
    .B(_1113_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_1 _3011_ (.A(net597),
    .B(_1115_),
    .Y(_0198_));
 sky130_fd_sc_hd__and4_1 _3012_ (.A(net278),
    .B(\scs.acc1[21] ),
    .C(_1110_),
    .D(_1112_),
    .X(_1116_));
 sky130_fd_sc_hd__xnor2_1 _3013_ (.A(net278),
    .B(_1114_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor2_1 _3014_ (.A(net597),
    .B(_1117_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _3015_ (.A(net277),
    .B(net60),
    .Y(_1118_));
 sky130_fd_sc_hd__xnor2_1 _3016_ (.A(net276),
    .B(net60),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_1 _3017_ (.A(net604),
    .B(_1119_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _3018_ (.A(_1468_),
    .B(_1118_),
    .Y(_1120_));
 sky130_fd_sc_hd__xnor2_1 _3019_ (.A(_1468_),
    .B(_1118_),
    .Y(_1121_));
 sky130_fd_sc_hd__nor2_1 _3020_ (.A(net604),
    .B(_1121_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand4_2 _3021_ (.A(net274),
    .B(net275),
    .C(net277),
    .D(net60),
    .Y(_1122_));
 sky130_fd_sc_hd__o211a_1 _3022_ (.A1(net274),
    .A2(_1120_),
    .B1(_1122_),
    .C1(net570),
    .X(_0202_));
 sky130_fd_sc_hd__xnor2_1 _3023_ (.A(_1467_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor2_1 _3024_ (.A(net601),
    .B(_1123_),
    .Y(_0203_));
 sky130_fd_sc_hd__o21ba_1 _3025_ (.A1(_1467_),
    .A2(_1122_),
    .B1_N(net860),
    .X(_1124_));
 sky130_fd_sc_hd__and4_1 _3026_ (.A(\scs.acc1[27] ),
    .B(\scs.acc1[26] ),
    .C(\scs.acc1[25] ),
    .D(net275),
    .X(_1125_));
 sky130_fd_sc_hd__and3_1 _3027_ (.A(net277),
    .B(net60),
    .C(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nor3_1 _3028_ (.A(net601),
    .B(_1124_),
    .C(_1126_),
    .Y(_0204_));
 sky130_fd_sc_hd__xnor2_1 _3029_ (.A(net660),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__nor2_1 _3030_ (.A(net601),
    .B(_1127_),
    .Y(_0205_));
 sky130_fd_sc_hd__a21oi_1 _3031_ (.A1(net273),
    .A2(_1126_),
    .B1(net737),
    .Y(_1128_));
 sky130_fd_sc_hd__and2_1 _3032_ (.A(\scs.acc1[29] ),
    .B(net273),
    .X(_1129_));
 sky130_fd_sc_hd__and4_1 _3033_ (.A(net277),
    .B(_1116_),
    .C(_1125_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__nor3_1 _3034_ (.A(net601),
    .B(_1128_),
    .C(_1130_),
    .Y(_0206_));
 sky130_fd_sc_hd__xnor2_1 _3035_ (.A(net272),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__nor2_1 _3036_ (.A(net602),
    .B(_1131_),
    .Y(_0207_));
 sky130_fd_sc_hd__a21oi_1 _3037_ (.A1(net272),
    .A2(_1130_),
    .B1(net655),
    .Y(_1132_));
 sky130_fd_sc_hd__and3_1 _3038_ (.A(net655),
    .B(\scs.acc1[30] ),
    .C(_1130_),
    .X(_1133_));
 sky130_fd_sc_hd__nor3_1 _3039_ (.A(net602),
    .B(_1132_),
    .C(_1133_),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2b_1 _3040_ (.A_N(\scs.diff2[0] ),
    .B(\scs.diff2_d[0] ),
    .Y(_1134_));
 sky130_fd_sc_hd__and2b_1 _3041_ (.A_N(\scs.diff2_d[0] ),
    .B(\scs.diff2[0] ),
    .X(_1135_));
 sky130_fd_sc_hd__or3b_1 _3042_ (.A(_1135_),
    .B(net71),
    .C_N(_1134_),
    .X(_1136_));
 sky130_fd_sc_hd__o211a_1 _3043_ (.A1(net633),
    .A2(net149),
    .B1(_1136_),
    .C1(net473),
    .X(_0209_));
 sky130_fd_sc_hd__and2b_1 _3044_ (.A_N(\scs.diff2_d[1] ),
    .B(\scs.diff2[1] ),
    .X(_1137_));
 sky130_fd_sc_hd__nand2b_1 _3045_ (.A_N(\scs.diff2[1] ),
    .B(\scs.diff2_d[1] ),
    .Y(_1138_));
 sky130_fd_sc_hd__and2b_1 _3046_ (.A_N(_1137_),
    .B(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__xnor2_1 _3047_ (.A(_1134_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _3048_ (.A(net149),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__o211a_1 _3049_ (.A1(net632),
    .A2(net149),
    .B1(_1141_),
    .C1(net473),
    .X(_0210_));
 sky130_fd_sc_hd__nand2b_1 _3050_ (.A_N(\scs.diff2[2] ),
    .B(\scs.diff2_d[2] ),
    .Y(_1142_));
 sky130_fd_sc_hd__inv_2 _3051_ (.A(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2b_1 _3052_ (.A_N(\scs.diff2_d[2] ),
    .B(\scs.diff2[2] ),
    .Y(_1144_));
 sky130_fd_sc_hd__a21oi_2 _3053_ (.A1(_1134_),
    .A2(_1138_),
    .B1(_1137_),
    .Y(_1145_));
 sky130_fd_sc_hd__a21oi_1 _3054_ (.A1(_1142_),
    .A2(_1144_),
    .B1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__a31o_1 _3055_ (.A1(_1142_),
    .A2(_1144_),
    .A3(_1145_),
    .B1(net72),
    .X(_1147_));
 sky130_fd_sc_hd__o221a_1 _3056_ (.A1(net664),
    .A2(net152),
    .B1(_1146_),
    .B2(_1147_),
    .C1(net473),
    .X(_0211_));
 sky130_fd_sc_hd__o21ai_2 _3057_ (.A1(_1143_),
    .A2(_1145_),
    .B1(_1144_),
    .Y(_1148_));
 sky130_fd_sc_hd__nand2b_1 _3058_ (.A_N(\scs.diff2[3] ),
    .B(\scs.diff2_d[3] ),
    .Y(_1149_));
 sky130_fd_sc_hd__inv_2 _3059_ (.A(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__and2b_1 _3060_ (.A_N(\scs.diff2_d[3] ),
    .B(\scs.diff2[3] ),
    .X(_1151_));
 sky130_fd_sc_hd__o21a_1 _3061_ (.A1(_1150_),
    .A2(_1151_),
    .B1(_1148_),
    .X(_1152_));
 sky130_fd_sc_hd__o31ai_1 _3062_ (.A1(_1148_),
    .A2(_1150_),
    .A3(_1151_),
    .B1(net150),
    .Y(_1153_));
 sky130_fd_sc_hd__o221a_1 _3063_ (.A1(net644),
    .A2(net150),
    .B1(_1152_),
    .B2(_1153_),
    .C1(net474),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_1 _3064_ (.A1(_1148_),
    .A2(_1149_),
    .B1(_1151_),
    .X(_1154_));
 sky130_fd_sc_hd__and2b_1 _3065_ (.A_N(\scs.diff2_d[4] ),
    .B(\scs.diff2[4] ),
    .X(_1155_));
 sky130_fd_sc_hd__and2b_1 _3066_ (.A_N(\scs.diff2[4] ),
    .B(\scs.diff2_d[4] ),
    .X(_1156_));
 sky130_fd_sc_hd__nor2_1 _3067_ (.A(_1155_),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__xor2_1 _3068_ (.A(_1154_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__or2_1 _3069_ (.A(net758),
    .B(net150),
    .X(_1159_));
 sky130_fd_sc_hd__o211a_1 _3070_ (.A1(net72),
    .A2(_1158_),
    .B1(_1159_),
    .C1(net478),
    .X(_0213_));
 sky130_fd_sc_hd__nand2b_1 _3071_ (.A_N(\scs.diff2[5] ),
    .B(\scs.diff2_d[5] ),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2b_1 _3072_ (.A_N(\scs.diff2_d[5] ),
    .B(\scs.diff2[5] ),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _3073_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__a21o_1 _3075_ (.A1(_1154_),
    .A2(_1157_),
    .B1(_1155_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_1 _3076_ (.A(_1162_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21o_1 _3077_ (.A1(_1162_),
    .A2(_1164_),
    .B1(net73),
    .X(_1166_));
 sky130_fd_sc_hd__o221a_1 _3078_ (.A1(net646),
    .A2(net156),
    .B1(_1165_),
    .B2(_1166_),
    .C1(net478),
    .X(_0214_));
 sky130_fd_sc_hd__a21bo_1 _3079_ (.A1(_1155_),
    .A2(_1160_),
    .B1_N(_1161_),
    .X(_1167_));
 sky130_fd_sc_hd__a31o_1 _3080_ (.A1(_1154_),
    .A2(_1157_),
    .A3(_1163_),
    .B1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__and2b_1 _3081_ (.A_N(\scs.diff2_d[6] ),
    .B(\scs.diff2[6] ),
    .X(_1169_));
 sky130_fd_sc_hd__and2b_1 _3082_ (.A_N(\scs.diff2[6] ),
    .B(\scs.diff2_d[6] ),
    .X(_1170_));
 sky130_fd_sc_hd__nor2_1 _3083_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _3084_ (.A(_1168_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(_1168_),
    .B(_1171_),
    .X(_1173_));
 sky130_fd_sc_hd__a21o_1 _3086_ (.A1(_1172_),
    .A2(_1173_),
    .B1(net75),
    .X(_1174_));
 sky130_fd_sc_hd__o211a_1 _3087_ (.A1(net631),
    .A2(net156),
    .B1(_1174_),
    .C1(net479),
    .X(_0215_));
 sky130_fd_sc_hd__nand2b_1 _3088_ (.A_N(net424),
    .B(\scs.diff2_d[7] ),
    .Y(_1175_));
 sky130_fd_sc_hd__and2b_1 _3089_ (.A_N(\scs.diff2_d[7] ),
    .B(net424),
    .X(_1176_));
 sky130_fd_sc_hd__nand2b_1 _3090_ (.A_N(\scs.diff2_d[7] ),
    .B(net424),
    .Y(_1177_));
 sky130_fd_sc_hd__nand2_1 _3091_ (.A(_1175_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__a21o_1 _3092_ (.A1(_1168_),
    .A2(_1171_),
    .B1(_1169_),
    .X(_1179_));
 sky130_fd_sc_hd__nor2_1 _3093_ (.A(_1178_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__a21o_1 _3094_ (.A1(_1178_),
    .A2(_1179_),
    .B1(net76),
    .X(_1181_));
 sky130_fd_sc_hd__o221a_1 _3095_ (.A1(net642),
    .A2(net156),
    .B1(_1180_),
    .B2(_1181_),
    .C1(net479),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _3096_ (.A(_1169_),
    .B(_1175_),
    .X(_1182_));
 sky130_fd_sc_hd__a311o_1 _3097_ (.A1(_1168_),
    .A2(_1171_),
    .A3(_1175_),
    .B1(_1176_),
    .C1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__and2b_1 _3098_ (.A_N(\scs.diff2_d[8] ),
    .B(\scs.diff2[8] ),
    .X(_1184_));
 sky130_fd_sc_hd__and2b_1 _3099_ (.A_N(\scs.diff2[8] ),
    .B(\scs.diff2_d[8] ),
    .X(_1185_));
 sky130_fd_sc_hd__nor2_1 _3100_ (.A(_1184_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__xor2_1 _3101_ (.A(_1183_),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__or2_1 _3102_ (.A(net749),
    .B(net171),
    .X(_1188_));
 sky130_fd_sc_hd__o211a_1 _3103_ (.A1(net75),
    .A2(_1187_),
    .B1(_1188_),
    .C1(net491),
    .X(_0217_));
 sky130_fd_sc_hd__nand2b_2 _3104_ (.A_N(\scs.diff2[9] ),
    .B(\scs.diff2_d[9] ),
    .Y(_1189_));
 sky130_fd_sc_hd__inv_2 _3105_ (.A(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__and2b_1 _3106_ (.A_N(\scs.diff2_d[9] ),
    .B(\scs.diff2[9] ),
    .X(_1191_));
 sky130_fd_sc_hd__nor2_1 _3107_ (.A(_1190_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__a21oi_1 _3108_ (.A1(_1183_),
    .A2(_1186_),
    .B1(_1184_),
    .Y(_1193_));
 sky130_fd_sc_hd__and2_1 _3109_ (.A(_1192_),
    .B(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__o21ai_1 _3110_ (.A1(_1192_),
    .A2(_1193_),
    .B1(net171),
    .Y(_1195_));
 sky130_fd_sc_hd__o221a_1 _3111_ (.A1(net641),
    .A2(net171),
    .B1(_1194_),
    .B2(_1195_),
    .C1(net491),
    .X(_0218_));
 sky130_fd_sc_hd__nand2b_1 _3112_ (.A_N(\scs.diff2_d[10] ),
    .B(\scs.diff2[10] ),
    .Y(_1196_));
 sky130_fd_sc_hd__inv_2 _3113_ (.A(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2b_1 _3114_ (.A_N(\scs.diff2[10] ),
    .B(\scs.diff2_d[10] ),
    .Y(_1198_));
 sky130_fd_sc_hd__a211o_1 _3115_ (.A1(_1183_),
    .A2(_1186_),
    .B1(_1191_),
    .C1(_1184_),
    .X(_1199_));
 sky130_fd_sc_hd__a22oi_1 _3116_ (.A1(_1196_),
    .A2(_1198_),
    .B1(_1199_),
    .B2(_1189_),
    .Y(_1200_));
 sky130_fd_sc_hd__a41o_1 _3117_ (.A1(_1189_),
    .A2(_1196_),
    .A3(_1198_),
    .A4(_1199_),
    .B1(net89),
    .X(_1201_));
 sky130_fd_sc_hd__o2bb2a_1 _3118_ (.A1_N(net852),
    .A2_N(net88),
    .B1(_1200_),
    .B2(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__nor2_1 _3119_ (.A(net592),
    .B(_1202_),
    .Y(_0219_));
 sky130_fd_sc_hd__and2b_1 _3120_ (.A_N(\scs.diff2_d[11] ),
    .B(\scs.diff2[11] ),
    .X(_1203_));
 sky130_fd_sc_hd__nand2b_1 _3121_ (.A_N(\scs.diff2[11] ),
    .B(\scs.diff2_d[11] ),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2b_1 _3122_ (.A_N(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__a31o_1 _3123_ (.A1(_1189_),
    .A2(_1198_),
    .A3(_1199_),
    .B1(_1197_),
    .X(_1206_));
 sky130_fd_sc_hd__xnor2_1 _3124_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(net800),
    .A1(_1207_),
    .S(net172),
    .X(_1208_));
 sky130_fd_sc_hd__and2_1 _3126_ (.A(net491),
    .B(_1208_),
    .X(_0220_));
 sky130_fd_sc_hd__a21oi_2 _3127_ (.A1(_1204_),
    .A2(_1206_),
    .B1(_1203_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2b_1 _3128_ (.A_N(\scs.diff2_d[12] ),
    .B(\scs.diff2[12] ),
    .Y(_1210_));
 sky130_fd_sc_hd__nand2b_1 _3129_ (.A_N(\scs.diff2[12] ),
    .B(\scs.diff2_d[12] ),
    .Y(_1211_));
 sky130_fd_sc_hd__nand2_1 _3130_ (.A(_1210_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__or2_1 _3131_ (.A(_1209_),
    .B(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__xnor2_1 _3132_ (.A(_1209_),
    .B(_1212_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _3133_ (.A(net176),
    .B(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__o211a_1 _3134_ (.A1(net628),
    .A2(net176),
    .B1(_1215_),
    .C1(net495),
    .X(_0221_));
 sky130_fd_sc_hd__and2b_1 _3135_ (.A_N(\scs.diff2[13] ),
    .B(\scs.diff2_d[13] ),
    .X(_1216_));
 sky130_fd_sc_hd__nand2b_1 _3136_ (.A_N(\scs.diff2_d[13] ),
    .B(\scs.diff2[13] ),
    .Y(_1217_));
 sky130_fd_sc_hd__and2b_1 _3137_ (.A_N(_1216_),
    .B(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__inv_2 _3138_ (.A(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__a21oi_1 _3139_ (.A1(_1210_),
    .A2(_1213_),
    .B1(_1218_),
    .Y(_1220_));
 sky130_fd_sc_hd__a31o_1 _3140_ (.A1(_1210_),
    .A2(_1213_),
    .A3(_1218_),
    .B1(net93),
    .X(_1221_));
 sky130_fd_sc_hd__o221a_1 _3141_ (.A1(net643),
    .A2(net176),
    .B1(_1220_),
    .B2(_1221_),
    .C1(net495),
    .X(_0222_));
 sky130_fd_sc_hd__nand2b_1 _3142_ (.A_N(\scs.diff2_d[14] ),
    .B(\scs.diff2[14] ),
    .Y(_1222_));
 sky130_fd_sc_hd__nand2b_1 _3143_ (.A_N(\scs.diff2[14] ),
    .B(\scs.diff2_d[14] ),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _3144_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__or2_1 _3145_ (.A(_1210_),
    .B(_1216_),
    .X(_1225_));
 sky130_fd_sc_hd__o311a_1 _3146_ (.A1(_1209_),
    .A2(_1212_),
    .A3(_1219_),
    .B1(_1225_),
    .C1(_1217_),
    .X(_1226_));
 sky130_fd_sc_hd__or2_1 _3147_ (.A(_1224_),
    .B(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__xor2_1 _3148_ (.A(_1224_),
    .B(_1226_),
    .X(_1228_));
 sky130_fd_sc_hd__or2_1 _3149_ (.A(net767),
    .B(net177),
    .X(_1229_));
 sky130_fd_sc_hd__o211a_1 _3150_ (.A1(net92),
    .A2(_1228_),
    .B1(_1229_),
    .C1(net495),
    .X(_0223_));
 sky130_fd_sc_hd__xnor2_1 _3151_ (.A(\scs.diff2_d[15] ),
    .B(net423),
    .Y(_1230_));
 sky130_fd_sc_hd__inv_2 _3152_ (.A(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__a21oi_1 _3153_ (.A1(_1222_),
    .A2(_1227_),
    .B1(_1230_),
    .Y(_1232_));
 sky130_fd_sc_hd__a31o_1 _3154_ (.A1(_1222_),
    .A2(_1227_),
    .A3(_1230_),
    .B1(net92),
    .X(_1233_));
 sky130_fd_sc_hd__o221a_1 _3155_ (.A1(net645),
    .A2(net180),
    .B1(_1232_),
    .B2(_1233_),
    .C1(net496),
    .X(_0224_));
 sky130_fd_sc_hd__nand2b_1 _3156_ (.A_N(\scs.diff2_d[16] ),
    .B(\scs.diff2[16] ),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2b_1 _3157_ (.A_N(\scs.diff2[16] ),
    .B(\scs.diff2_d[16] ),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _3158_ (.A(_1234_),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__o21ba_1 _3159_ (.A1(_1460_),
    .A2(net423),
    .B1_N(_1222_),
    .X(_1237_));
 sky130_fd_sc_hd__a21oi_1 _3160_ (.A1(_1460_),
    .A2(net423),
    .B1(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__o31a_1 _3161_ (.A1(_1224_),
    .A2(_1226_),
    .A3(_1231_),
    .B1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__or2_1 _3162_ (.A(_1236_),
    .B(net64),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _3163_ (.A(_1236_),
    .B(net64),
    .Y(_1241_));
 sky130_fd_sc_hd__a21o_1 _3164_ (.A1(_1240_),
    .A2(_1241_),
    .B1(net109),
    .X(_1242_));
 sky130_fd_sc_hd__o211a_1 _3165_ (.A1(net630),
    .A2(net193),
    .B1(_1242_),
    .C1(net522),
    .X(_0225_));
 sky130_fd_sc_hd__and2b_1 _3166_ (.A_N(\scs.diff2_d[17] ),
    .B(net422),
    .X(_1243_));
 sky130_fd_sc_hd__nand2b_1 _3167_ (.A_N(\scs.diff2_d[17] ),
    .B(net422),
    .Y(_1244_));
 sky130_fd_sc_hd__and2b_1 _3168_ (.A_N(net422),
    .B(\scs.diff2_d[17] ),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_1 _3169_ (.A(_1243_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__o21a_1 _3170_ (.A1(_1236_),
    .A2(net64),
    .B1(_1234_),
    .X(_1247_));
 sky130_fd_sc_hd__xnor2_1 _3171_ (.A(_1246_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__or2_1 _3172_ (.A(net746),
    .B(net193),
    .X(_1249_));
 sky130_fd_sc_hd__o211a_1 _3173_ (.A1(net109),
    .A2(_1248_),
    .B1(_1249_),
    .C1(net523),
    .X(_0226_));
 sky130_fd_sc_hd__nand2b_1 _3174_ (.A_N(\scs.diff2_d[18] ),
    .B(net421),
    .Y(_1250_));
 sky130_fd_sc_hd__xnor2_2 _3175_ (.A(\scs.diff2_d[18] ),
    .B(net421),
    .Y(_1251_));
 sky130_fd_sc_hd__inv_2 _3176_ (.A(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21o_1 _3177_ (.A1(_1244_),
    .A2(_1247_),
    .B1(_1245_),
    .X(_1253_));
 sky130_fd_sc_hd__or2_1 _3178_ (.A(_1252_),
    .B(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__xnor2_1 _3179_ (.A(_1251_),
    .B(_1253_),
    .Y(_1255_));
 sky130_fd_sc_hd__or2_1 _3180_ (.A(net748),
    .B(net194),
    .X(_1256_));
 sky130_fd_sc_hd__o211a_1 _3181_ (.A1(net108),
    .A2(_1255_),
    .B1(_1256_),
    .C1(net522),
    .X(_0227_));
 sky130_fd_sc_hd__xnor2_1 _3182_ (.A(\scs.diff2_d[19] ),
    .B(net420),
    .Y(_1257_));
 sky130_fd_sc_hd__a21oi_1 _3183_ (.A1(_1250_),
    .A2(_1254_),
    .B1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__a31o_1 _3184_ (.A1(_1250_),
    .A2(_1254_),
    .A3(_1257_),
    .B1(net108),
    .X(_1259_));
 sky130_fd_sc_hd__o221a_1 _3185_ (.A1(net635),
    .A2(net193),
    .B1(_1258_),
    .B2(_1259_),
    .C1(net523),
    .X(_0228_));
 sky130_fd_sc_hd__and2b_1 _3186_ (.A_N(\scs.diff2_d[20] ),
    .B(\scs.diff2[20] ),
    .X(_1260_));
 sky130_fd_sc_hd__and2b_1 _3187_ (.A_N(\scs.diff2[20] ),
    .B(\scs.diff2_d[20] ),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_1 _3188_ (.A(_1260_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _3189_ (.A(_1251_),
    .B(_1257_),
    .Y(_1263_));
 sky130_fd_sc_hd__a211o_1 _3190_ (.A1(_1234_),
    .A2(_1244_),
    .B1(_1245_),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__o21ai_1 _3191_ (.A1(_1458_),
    .A2(net420),
    .B1(net421),
    .Y(_1265_));
 sky130_fd_sc_hd__o221a_1 _3192_ (.A1(\scs.diff2_d[19] ),
    .A2(_1459_),
    .B1(\scs.diff2_d[18] ),
    .B2(_1265_),
    .C1(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__or4_1 _3193_ (.A(_1236_),
    .B(_1243_),
    .C(_1245_),
    .D(_1263_),
    .X(_1267_));
 sky130_fd_sc_hd__o21ai_1 _3194_ (.A1(_1239_),
    .A2(_1267_),
    .B1(_1266_),
    .Y(_1268_));
 sky130_fd_sc_hd__xnor2_1 _3195_ (.A(_1262_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__nor2_1 _3196_ (.A(net701),
    .B(net197),
    .Y(_1270_));
 sky130_fd_sc_hd__a211oi_1 _3197_ (.A1(net197),
    .A2(_1269_),
    .B1(_1270_),
    .C1(net593),
    .Y(_0229_));
 sky130_fd_sc_hd__and2b_1 _3198_ (.A_N(\scs.diff2_d[21] ),
    .B(net419),
    .X(_1271_));
 sky130_fd_sc_hd__nand2b_1 _3199_ (.A_N(\scs.diff2_d[21] ),
    .B(net419),
    .Y(_1272_));
 sky130_fd_sc_hd__and2b_1 _3200_ (.A_N(net419),
    .B(\scs.diff2_d[21] ),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(_1271_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__a21oi_1 _3202_ (.A1(_1262_),
    .A2(_1268_),
    .B1(_1260_),
    .Y(_1275_));
 sky130_fd_sc_hd__and2_1 _3203_ (.A(_1274_),
    .B(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__o21ai_1 _3204_ (.A1(_1274_),
    .A2(_1275_),
    .B1(net197),
    .Y(_1277_));
 sky130_fd_sc_hd__o221a_1 _3205_ (.A1(net634),
    .A2(net197),
    .B1(_1276_),
    .B2(_1277_),
    .C1(net528),
    .X(_0230_));
 sky130_fd_sc_hd__nand2b_1 _3206_ (.A_N(\scs.diff2_d[22] ),
    .B(\scs.diff2[22] ),
    .Y(_1278_));
 sky130_fd_sc_hd__nand2b_1 _3207_ (.A_N(\scs.diff2[22] ),
    .B(\scs.diff2_d[22] ),
    .Y(_1279_));
 sky130_fd_sc_hd__nand2_1 _3208_ (.A(_1278_),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__a21o_1 _3209_ (.A1(_1272_),
    .A2(_1275_),
    .B1(_1273_),
    .X(_1281_));
 sky130_fd_sc_hd__nand2_1 _3210_ (.A(_1280_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__or2_1 _3211_ (.A(_1280_),
    .B(_1281_),
    .X(_1283_));
 sky130_fd_sc_hd__a21o_1 _3212_ (.A1(_1282_),
    .A2(_1283_),
    .B1(net112),
    .X(_1284_));
 sky130_fd_sc_hd__o211a_1 _3213_ (.A1(net626),
    .A2(net198),
    .B1(_1284_),
    .C1(net528),
    .X(_0231_));
 sky130_fd_sc_hd__and2b_1 _3214_ (.A_N(\scs.diff2[23] ),
    .B(\scs.diff2_d[23] ),
    .X(_1285_));
 sky130_fd_sc_hd__nand2b_1 _3215_ (.A_N(\scs.diff2_d[23] ),
    .B(\scs.diff2[23] ),
    .Y(_1286_));
 sky130_fd_sc_hd__and2b_1 _3216_ (.A_N(_1285_),
    .B(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__a21oi_1 _3217_ (.A1(_1278_),
    .A2(_1283_),
    .B1(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__and3_1 _3218_ (.A(_1278_),
    .B(_1283_),
    .C(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__or2_1 _3219_ (.A(net747),
    .B(net213),
    .X(_1290_));
 sky130_fd_sc_hd__o311a_1 _3220_ (.A1(net112),
    .A2(_1288_),
    .A3(_1289_),
    .B1(_1290_),
    .C1(net536),
    .X(_0232_));
 sky130_fd_sc_hd__nand2b_1 _3221_ (.A_N(\scs.diff2_d[24] ),
    .B(\scs.diff2[24] ),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2b_1 _3222_ (.A_N(\scs.diff2[24] ),
    .B(\scs.diff2_d[24] ),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _3223_ (.A(_1291_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__nand2b_1 _3224_ (.A_N(_1280_),
    .B(_1287_),
    .Y(_1294_));
 sky130_fd_sc_hd__or4b_1 _3225_ (.A(_1271_),
    .B(_1273_),
    .C(_1294_),
    .D_N(_1262_),
    .X(_1295_));
 sky130_fd_sc_hd__nand2b_1 _3226_ (.A_N(_1273_),
    .B(_1260_),
    .Y(_1296_));
 sky130_fd_sc_hd__a21o_1 _3227_ (.A1(_1272_),
    .A2(_1296_),
    .B1(_1294_),
    .X(_1297_));
 sky130_fd_sc_hd__a21o_1 _3228_ (.A1(_1278_),
    .A2(_1286_),
    .B1(_1285_),
    .X(_1298_));
 sky130_fd_sc_hd__o211a_1 _3229_ (.A1(_1266_),
    .A2(_1295_),
    .B1(_1297_),
    .C1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o31a_1 _3230_ (.A1(net64),
    .A2(_1267_),
    .A3(_1295_),
    .B1(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__or2_1 _3231_ (.A(_1293_),
    .B(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _3232_ (.A(_1293_),
    .B(_1300_),
    .Y(_1302_));
 sky130_fd_sc_hd__a21o_1 _3233_ (.A1(_1301_),
    .A2(_1302_),
    .B1(net123),
    .X(_1303_));
 sky130_fd_sc_hd__o211a_1 _3234_ (.A1(net627),
    .A2(net213),
    .B1(_1303_),
    .C1(net536),
    .X(_0233_));
 sky130_fd_sc_hd__nand2b_1 _3235_ (.A_N(\scs.diff2_d[25] ),
    .B(\scs.diff2[25] ),
    .Y(_1304_));
 sky130_fd_sc_hd__and2b_1 _3236_ (.A_N(\scs.diff2[25] ),
    .B(\scs.diff2_d[25] ),
    .X(_1305_));
 sky130_fd_sc_hd__inv_2 _3237_ (.A(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _3238_ (.A(_1304_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__nand2_1 _3239_ (.A(_1291_),
    .B(_1301_),
    .Y(_1308_));
 sky130_fd_sc_hd__xnor2_1 _3240_ (.A(_1307_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__or2_1 _3241_ (.A(net759),
    .B(net213),
    .X(_1310_));
 sky130_fd_sc_hd__o211a_1 _3242_ (.A1(net123),
    .A2(_1309_),
    .B1(_1310_),
    .C1(net537),
    .X(_0234_));
 sky130_fd_sc_hd__nand2b_1 _3243_ (.A_N(\scs.diff2_d[26] ),
    .B(\scs.diff2[26] ),
    .Y(_1311_));
 sky130_fd_sc_hd__xnor2_2 _3244_ (.A(\scs.diff2_d[26] ),
    .B(\scs.diff2[26] ),
    .Y(_1312_));
 sky130_fd_sc_hd__inv_2 _3245_ (.A(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a31o_1 _3246_ (.A1(_1291_),
    .A2(_1301_),
    .A3(_1304_),
    .B1(_1305_),
    .X(_1314_));
 sky130_fd_sc_hd__or2_1 _3247_ (.A(_1313_),
    .B(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__xnor2_1 _3248_ (.A(_1312_),
    .B(_1314_),
    .Y(_1316_));
 sky130_fd_sc_hd__or2_1 _3249_ (.A(net752),
    .B(net214),
    .X(_1317_));
 sky130_fd_sc_hd__o211a_1 _3250_ (.A1(net124),
    .A2(_1316_),
    .B1(_1317_),
    .C1(net537),
    .X(_0235_));
 sky130_fd_sc_hd__xnor2_1 _3251_ (.A(\scs.diff2_d[27] ),
    .B(\scs.diff2[27] ),
    .Y(_1318_));
 sky130_fd_sc_hd__a21oi_1 _3252_ (.A1(_1311_),
    .A2(_1315_),
    .B1(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__a31o_1 _3253_ (.A1(_1311_),
    .A2(_1315_),
    .A3(_1318_),
    .B1(net129),
    .X(_1320_));
 sky130_fd_sc_hd__o221a_1 _3254_ (.A1(net647),
    .A2(net217),
    .B1(_1319_),
    .B2(_1320_),
    .C1(net537),
    .X(_0236_));
 sky130_fd_sc_hd__nand2_1 _3255_ (.A(_1312_),
    .B(_1318_),
    .Y(_1321_));
 sky130_fd_sc_hd__or4_1 _3256_ (.A(_1293_),
    .B(_1300_),
    .C(_1307_),
    .D(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a211o_1 _3257_ (.A1(_1291_),
    .A2(_1304_),
    .B1(_1305_),
    .C1(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__a21o_1 _3258_ (.A1(\scs.diff2_d[27] ),
    .A2(_1457_),
    .B1(_1311_),
    .X(_1324_));
 sky130_fd_sc_hd__o2111a_1 _3259_ (.A1(\scs.diff2_d[27] ),
    .A2(_1457_),
    .B1(_1322_),
    .C1(_1323_),
    .D1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__and2b_1 _3260_ (.A_N(\scs.diff2[28] ),
    .B(\scs.diff2_d[28] ),
    .X(_1326_));
 sky130_fd_sc_hd__nand2b_1 _3261_ (.A_N(\scs.diff2_d[28] ),
    .B(\scs.diff2[28] ),
    .Y(_1327_));
 sky130_fd_sc_hd__and2b_1 _3262_ (.A_N(_1326_),
    .B(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__and2_1 _3263_ (.A(_1325_),
    .B(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__o21ai_1 _3264_ (.A1(_1325_),
    .A2(_1328_),
    .B1(net217),
    .Y(_1330_));
 sky130_fd_sc_hd__o221a_1 _3265_ (.A1(net649),
    .A2(net217),
    .B1(_1329_),
    .B2(_1330_),
    .C1(net541),
    .X(_0237_));
 sky130_fd_sc_hd__o21ai_1 _3266_ (.A1(_1325_),
    .A2(_1326_),
    .B1(_1327_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2b_1 _3267_ (.A_N(\scs.diff2[29] ),
    .B(\scs.diff2_d[29] ),
    .Y(_1332_));
 sky130_fd_sc_hd__nand2b_1 _3268_ (.A_N(\scs.diff2_d[29] ),
    .B(\scs.diff2[29] ),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _3269_ (.A(_1332_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_1 _3270_ (.A(_1331_),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__a21o_1 _3271_ (.A1(_1331_),
    .A2(_1334_),
    .B1(net127),
    .X(_1336_));
 sky130_fd_sc_hd__o221a_1 _3272_ (.A1(net648),
    .A2(net218),
    .B1(_1335_),
    .B2(_1336_),
    .C1(net541),
    .X(_0238_));
 sky130_fd_sc_hd__nand2b_1 _3273_ (.A_N(\scs.diff2_d[30] ),
    .B(\scs.diff2[30] ),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2b_1 _3274_ (.A_N(\scs.diff2[30] ),
    .B(\scs.diff2_d[30] ),
    .Y(_1338_));
 sky130_fd_sc_hd__a21bo_1 _3275_ (.A1(_1331_),
    .A2(_1332_),
    .B1_N(_1333_),
    .X(_1339_));
 sky130_fd_sc_hd__a21o_1 _3276_ (.A1(_1337_),
    .A2(_1338_),
    .B1(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__a31oi_1 _3277_ (.A1(_1337_),
    .A2(_1338_),
    .A3(_1339_),
    .B1(net127),
    .Y(_1341_));
 sky130_fd_sc_hd__a22o_1 _3278_ (.A1(net813),
    .A2(net127),
    .B1(_1340_),
    .B2(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__and2_1 _3279_ (.A(net541),
    .B(_1342_),
    .X(_0239_));
 sky130_fd_sc_hd__a21bo_1 _3280_ (.A1(_1338_),
    .A2(_1339_),
    .B1_N(_1337_),
    .X(_1343_));
 sky130_fd_sc_hd__xor2_1 _3281_ (.A(\scs.diff2_d[31] ),
    .B(\scs.diff2[31] ),
    .X(_1344_));
 sky130_fd_sc_hd__xnor2_1 _3282_ (.A(_1343_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__or2_1 _3283_ (.A(net768),
    .B(net218),
    .X(_1346_));
 sky130_fd_sc_hd__o211a_1 _3284_ (.A1(net127),
    .A2(_1345_),
    .B1(_1346_),
    .C1(net542),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _3285_ (.A(net710),
    .B(net161),
    .X(_1347_));
 sky130_fd_sc_hd__o211a_1 _3286_ (.A1(net751),
    .A2(net81),
    .B1(_1347_),
    .C1(net484),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _3287_ (.A(\scs.diff1_d[1] ),
    .B(net161),
    .X(_1348_));
 sky130_fd_sc_hd__o211a_1 _3288_ (.A1(net693),
    .A2(net81),
    .B1(_1348_),
    .C1(net484),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _3289_ (.A(\scs.diff1_d[2] ),
    .B(net162),
    .X(_1349_));
 sky130_fd_sc_hd__o211a_1 _3290_ (.A1(net668),
    .A2(net81),
    .B1(_1349_),
    .C1(net485),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _3291_ (.A(\scs.diff1_d[3] ),
    .B(net154),
    .X(_1350_));
 sky130_fd_sc_hd__o211a_1 _3292_ (.A1(net678),
    .A2(net73),
    .B1(_1350_),
    .C1(net485),
    .X(_0244_));
 sky130_fd_sc_hd__or2_1 _3293_ (.A(\scs.diff1_d[4] ),
    .B(net166),
    .X(_1351_));
 sky130_fd_sc_hd__o211a_1 _3294_ (.A1(net702),
    .A2(net82),
    .B1(_1351_),
    .C1(net485),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _3295_ (.A(\scs.diff1_d[5] ),
    .B(net166),
    .X(_1352_));
 sky130_fd_sc_hd__o211a_1 _3296_ (.A1(net742),
    .A2(net82),
    .B1(_1352_),
    .C1(net486),
    .X(_0246_));
 sky130_fd_sc_hd__or2_1 _3297_ (.A(\scs.diff1_d[6] ),
    .B(net167),
    .X(_1353_));
 sky130_fd_sc_hd__o211a_1 _3298_ (.A1(net704),
    .A2(net83),
    .B1(_1353_),
    .C1(net486),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _3299_ (.A(net827),
    .B(net158),
    .X(_1354_));
 sky130_fd_sc_hd__o211a_1 _3300_ (.A1(net418),
    .A2(net77),
    .B1(_1354_),
    .C1(net494),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _3301_ (.A(\scs.diff1_d[8] ),
    .B(net182),
    .X(_1355_));
 sky130_fd_sc_hd__o211a_1 _3302_ (.A1(net676),
    .A2(net98),
    .B1(_1355_),
    .C1(net500),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _3303_ (.A(\scs.diff1_d[9] ),
    .B(net173),
    .X(_1356_));
 sky130_fd_sc_hd__o211a_1 _3304_ (.A1(net670),
    .A2(net90),
    .B1(_1356_),
    .C1(net501),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _3305_ (.A(net730),
    .B(net183),
    .X(_1357_));
 sky130_fd_sc_hd__o211a_1 _3306_ (.A1(net690),
    .A2(net99),
    .B1(_1357_),
    .C1(net501),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _3307_ (.A(net715),
    .B(net174),
    .X(_1358_));
 sky130_fd_sc_hd__o211a_1 _3308_ (.A1(net653),
    .A2(net90),
    .B1(_1358_),
    .C1(net497),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _3309_ (.A(\scs.diff1_d[12] ),
    .B(net186),
    .X(_1359_));
 sky130_fd_sc_hd__o211a_1 _3310_ (.A1(net716),
    .A2(net102),
    .B1(_1359_),
    .C1(net504),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _3311_ (.A(\scs.diff1_d[13] ),
    .B(net178),
    .X(_1360_));
 sky130_fd_sc_hd__o211a_1 _3312_ (.A1(net772),
    .A2(net94),
    .B1(_1360_),
    .C1(net504),
    .X(_0254_));
 sky130_fd_sc_hd__or2_1 _3313_ (.A(\scs.diff1_d[14] ),
    .B(net187),
    .X(_1361_));
 sky130_fd_sc_hd__o211a_1 _3314_ (.A1(net731),
    .A2(net103),
    .B1(_1361_),
    .C1(net530),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _3315_ (.A(_1466_),
    .B(net95),
    .Y(_1362_));
 sky130_fd_sc_hd__o211a_1 _3316_ (.A1(net417),
    .A2(net94),
    .B1(_1362_),
    .C1(net530),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _3317_ (.A(\scs.diff1_d[16] ),
    .B(net203),
    .X(_1363_));
 sky130_fd_sc_hd__o211a_1 _3318_ (.A1(net682),
    .A2(net115),
    .B1(_1363_),
    .C1(net530),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _3319_ (.A(net820),
    .B(net203),
    .X(_1364_));
 sky130_fd_sc_hd__o211a_1 _3320_ (.A1(net416),
    .A2(net115),
    .B1(_1364_),
    .C1(net530),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _3321_ (.A(\scs.diff1_d[18] ),
    .B(net204),
    .X(_1365_));
 sky130_fd_sc_hd__o211a_1 _3322_ (.A1(net415),
    .A2(net116),
    .B1(_1365_),
    .C1(net532),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _3323_ (.A(_1464_),
    .B(net116),
    .Y(_1366_));
 sky130_fd_sc_hd__o211a_1 _3324_ (.A1(net414),
    .A2(net116),
    .B1(_1366_),
    .C1(net532),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _3325_ (.A(\scs.diff1_d[20] ),
    .B(net208),
    .X(_1367_));
 sky130_fd_sc_hd__o211a_1 _3326_ (.A1(net665),
    .A2(net119),
    .B1(_1367_),
    .C1(net532),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _3327_ (.A(net817),
    .B(net207),
    .X(_1368_));
 sky130_fd_sc_hd__o211a_1 _3328_ (.A1(net413),
    .A2(net119),
    .B1(_1368_),
    .C1(net532),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _3329_ (.A(\scs.diff1_d[22] ),
    .B(net223),
    .X(_1369_));
 sky130_fd_sc_hd__o211a_1 _3330_ (.A1(net753),
    .A2(net134),
    .B1(_1369_),
    .C1(net548),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _3331_ (.A(net663),
    .B(net207),
    .X(_1370_));
 sky130_fd_sc_hd__o211a_1 _3332_ (.A1(net659),
    .A2(net134),
    .B1(_1370_),
    .C1(net548),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _3333_ (.A(\scs.diff1_d[24] ),
    .B(net223),
    .X(_1371_));
 sky130_fd_sc_hd__o211a_1 _3334_ (.A1(net686),
    .A2(net134),
    .B1(_1371_),
    .C1(net548),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _3335_ (.A(\scs.diff1_d[25] ),
    .B(net224),
    .X(_1372_));
 sky130_fd_sc_hd__o211a_1 _3336_ (.A1(net688),
    .A2(net135),
    .B1(_1372_),
    .C1(net548),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _3337_ (.A(\scs.diff1_d[26] ),
    .B(net227),
    .X(_1373_));
 sky130_fd_sc_hd__o211a_1 _3338_ (.A1(net835),
    .A2(net139),
    .B1(_1373_),
    .C1(net550),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _3339_ (.A(_1461_),
    .B(net139),
    .Y(_1374_));
 sky130_fd_sc_hd__o211a_1 _3340_ (.A1(\scs.diff1[27] ),
    .A2(net139),
    .B1(_1374_),
    .C1(net550),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _3341_ (.A(\scs.diff1_d[28] ),
    .B(net219),
    .X(_1375_));
 sky130_fd_sc_hd__o211a_1 _3342_ (.A1(net765),
    .A2(net131),
    .B1(_1375_),
    .C1(net550),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _3343_ (.A(\scs.diff1_d[29] ),
    .B(net228),
    .X(_1376_));
 sky130_fd_sc_hd__o211a_1 _3344_ (.A1(net726),
    .A2(net138),
    .B1(_1376_),
    .C1(net551),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _3345_ (.A(\scs.diff1_d[30] ),
    .B(net228),
    .X(_1377_));
 sky130_fd_sc_hd__o211a_1 _3346_ (.A1(net720),
    .A2(net138),
    .B1(_1377_),
    .C1(net551),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _3347_ (.A(\scs.diff1_d[31] ),
    .B(net228),
    .X(_1378_));
 sky130_fd_sc_hd__o211a_1 _3348_ (.A1(net661),
    .A2(net140),
    .B1(_1378_),
    .C1(net553),
    .X(_0272_));
 sky130_fd_sc_hd__or2_1 _3349_ (.A(net769),
    .B(net149),
    .X(_1379_));
 sky130_fd_sc_hd__o211a_1 _3350_ (.A1(net750),
    .A2(net71),
    .B1(_1379_),
    .C1(net473),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _3351_ (.A(\scs.diff2_d[1] ),
    .B(net153),
    .X(_1380_));
 sky130_fd_sc_hd__o211a_1 _3352_ (.A1(net699),
    .A2(net74),
    .B1(_1380_),
    .C1(net475),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _3353_ (.A(\scs.diff2_d[2] ),
    .B(net151),
    .X(_1381_));
 sky130_fd_sc_hd__o211a_1 _3354_ (.A1(net735),
    .A2(net71),
    .B1(_1381_),
    .C1(net476),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _3355_ (.A(\scs.diff2_d[3] ),
    .B(net150),
    .X(_1382_));
 sky130_fd_sc_hd__o211a_1 _3356_ (.A1(net756),
    .A2(net71),
    .B1(_1382_),
    .C1(net474),
    .X(_0276_));
 sky130_fd_sc_hd__or2_1 _3357_ (.A(\scs.diff2_d[4] ),
    .B(net151),
    .X(_1383_));
 sky130_fd_sc_hd__o211a_1 _3358_ (.A1(net672),
    .A2(net72),
    .B1(_1383_),
    .C1(net478),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _3359_ (.A(\scs.diff2_d[5] ),
    .B(net156),
    .X(_1384_));
 sky130_fd_sc_hd__o211a_1 _3360_ (.A1(net722),
    .A2(net75),
    .B1(_1384_),
    .C1(net478),
    .X(_0278_));
 sky130_fd_sc_hd__or2_1 _3361_ (.A(\scs.diff2_d[6] ),
    .B(net157),
    .X(_1385_));
 sky130_fd_sc_hd__o211a_1 _3362_ (.A1(net697),
    .A2(net76),
    .B1(_1385_),
    .C1(net479),
    .X(_0279_));
 sky130_fd_sc_hd__or2_1 _3363_ (.A(net828),
    .B(net157),
    .X(_1386_));
 sky130_fd_sc_hd__o211a_1 _3364_ (.A1(net424),
    .A2(net75),
    .B1(_1386_),
    .C1(net479),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _3365_ (.A(\scs.diff2_d[8] ),
    .B(net171),
    .X(_1387_));
 sky130_fd_sc_hd__o211a_1 _3366_ (.A1(net680),
    .A2(net88),
    .B1(_1387_),
    .C1(net491),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _3367_ (.A(\scs.diff2_d[9] ),
    .B(net172),
    .X(_1388_));
 sky130_fd_sc_hd__o211a_1 _3368_ (.A1(net728),
    .A2(net88),
    .B1(_1388_),
    .C1(net492),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _3369_ (.A(\scs.diff2_d[10] ),
    .B(net172),
    .X(_1389_));
 sky130_fd_sc_hd__o211a_1 _3370_ (.A1(net691),
    .A2(net88),
    .B1(_1389_),
    .C1(net492),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _3371_ (.A(\scs.diff2_d[11] ),
    .B(net175),
    .X(_1390_));
 sky130_fd_sc_hd__o211a_1 _3372_ (.A1(net674),
    .A2(net89),
    .B1(_1390_),
    .C1(net495),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(net739),
    .B(net177),
    .X(_1391_));
 sky130_fd_sc_hd__o211a_1 _3374_ (.A1(net733),
    .A2(net93),
    .B1(_1391_),
    .C1(net496),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _3375_ (.A(\scs.diff2_d[13] ),
    .B(net176),
    .X(_1392_));
 sky130_fd_sc_hd__o211a_1 _3376_ (.A1(net763),
    .A2(net93),
    .B1(_1392_),
    .C1(net496),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _3377_ (.A(\scs.diff2_d[14] ),
    .B(net177),
    .X(_1393_));
 sky130_fd_sc_hd__o211a_1 _3378_ (.A1(net621),
    .A2(net92),
    .B1(_1393_),
    .C1(net524),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _3379_ (.A(_1460_),
    .B(net92),
    .Y(_1394_));
 sky130_fd_sc_hd__o211a_1 _3380_ (.A1(net423),
    .A2(net96),
    .B1(_1394_),
    .C1(net522),
    .X(_0288_));
 sky130_fd_sc_hd__or2_1 _3381_ (.A(\scs.diff2_d[16] ),
    .B(net195),
    .X(_1395_));
 sky130_fd_sc_hd__o211a_1 _3382_ (.A1(net724),
    .A2(net110),
    .B1(_1395_),
    .C1(net525),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _3383_ (.A(net824),
    .B(net193),
    .X(_1396_));
 sky130_fd_sc_hd__o211a_1 _3384_ (.A1(net422),
    .A2(net109),
    .B1(_1396_),
    .C1(net522),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _3385_ (.A(\scs.diff2_d[18] ),
    .B(net194),
    .X(_1397_));
 sky130_fd_sc_hd__o211a_1 _3386_ (.A1(net421),
    .A2(net108),
    .B1(_1397_),
    .C1(net528),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _3387_ (.A(_1458_),
    .B(net108),
    .Y(_1398_));
 sky130_fd_sc_hd__o211a_1 _3388_ (.A1(net420),
    .A2(net111),
    .B1(_1398_),
    .C1(net527),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _3389_ (.A(\scs.diff2_d[20] ),
    .B(net199),
    .X(_1399_));
 sky130_fd_sc_hd__o211a_1 _3390_ (.A1(net718),
    .A2(net112),
    .B1(_1399_),
    .C1(net527),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _3391_ (.A(net815),
    .B(net198),
    .X(_1400_));
 sky130_fd_sc_hd__o211a_1 _3392_ (.A1(net419),
    .A2(net112),
    .B1(_1400_),
    .C1(net529),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _3393_ (.A(\scs.diff2_d[22] ),
    .B(net198),
    .X(_1401_));
 sky130_fd_sc_hd__o211a_1 _3394_ (.A1(net785),
    .A2(net123),
    .B1(_1401_),
    .C1(net536),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _3395_ (.A(\scs.diff2_d[23] ),
    .B(net200),
    .X(_1402_));
 sky130_fd_sc_hd__o211a_1 _3396_ (.A1(net684),
    .A2(net113),
    .B1(_1402_),
    .C1(net538),
    .X(_0296_));
 sky130_fd_sc_hd__or2_1 _3397_ (.A(net741),
    .B(net213),
    .X(_1403_));
 sky130_fd_sc_hd__o211a_1 _3398_ (.A1(net740),
    .A2(net123),
    .B1(_1403_),
    .C1(net536),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _3399_ (.A(\scs.diff2_d[25] ),
    .B(net214),
    .X(_1404_));
 sky130_fd_sc_hd__o211a_1 _3400_ (.A1(net713),
    .A2(net124),
    .B1(_1404_),
    .C1(net539),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _3401_ (.A(\scs.diff2_d[26] ),
    .B(net214),
    .X(_1405_));
 sky130_fd_sc_hd__o211a_1 _3402_ (.A1(net831),
    .A2(net124),
    .B1(_1405_),
    .C1(net539),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(_1456_),
    .B(net129),
    .Y(_1406_));
 sky130_fd_sc_hd__o211a_1 _3404_ (.A1(net846),
    .A2(net129),
    .B1(_1406_),
    .C1(net541),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _3405_ (.A(\scs.diff2_d[28] ),
    .B(net217),
    .X(_1407_));
 sky130_fd_sc_hd__o211a_1 _3406_ (.A1(net744),
    .A2(net129),
    .B1(_1407_),
    .C1(net543),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _3407_ (.A(\scs.diff2_d[29] ),
    .B(net218),
    .X(_1408_));
 sky130_fd_sc_hd__o211a_1 _3408_ (.A1(net783),
    .A2(net128),
    .B1(_1408_),
    .C1(net544),
    .X(_0302_));
 sky130_fd_sc_hd__or2_1 _3409_ (.A(\scs.diff2_d[30] ),
    .B(net218),
    .X(_1409_));
 sky130_fd_sc_hd__o211a_1 _3410_ (.A1(net777),
    .A2(net128),
    .B1(_1409_),
    .C1(net542),
    .X(_0303_));
 sky130_fd_sc_hd__or2_1 _3411_ (.A(\scs.diff2_d[31] ),
    .B(net220),
    .X(_1410_));
 sky130_fd_sc_hd__o211a_1 _3412_ (.A1(net707),
    .A2(net131),
    .B1(_1410_),
    .C1(net544),
    .X(_0304_));
 sky130_fd_sc_hd__o22a_1 _3413_ (.A1(_1453_),
    .A2(\scs.oversample_in[2] ),
    .B1(_1484_),
    .B2(\scs.word_count[9] ),
    .X(_1411_));
 sky130_fd_sc_hd__o22a_1 _3414_ (.A1(net267),
    .A2(_1480_),
    .B1(\scs.oversample_in[8] ),
    .B2(_1449_),
    .X(_1412_));
 sky130_fd_sc_hd__o22a_1 _3415_ (.A1(_1454_),
    .A2(\scs.oversample_in[1] ),
    .B1(_1481_),
    .B2(net265),
    .X(_1413_));
 sky130_fd_sc_hd__and3_1 _3416_ (.A(_1411_),
    .B(_1412_),
    .C(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__o221a_1 _3417_ (.A1(net268),
    .A2(_1479_),
    .B1(\scs.oversample_in[9] ),
    .B2(_1447_),
    .C1(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__xnor2_1 _3418_ (.A(net258),
    .B(\scs.oversample_in[6] ),
    .Y(_1416_));
 sky130_fd_sc_hd__xnor2_1 _3419_ (.A(net260),
    .B(\scs.oversample_in[5] ),
    .Y(_1417_));
 sky130_fd_sc_hd__xnor2_1 _3420_ (.A(net257),
    .B(\scs.oversample_in[7] ),
    .Y(_1418_));
 sky130_fd_sc_hd__xnor2_1 _3421_ (.A(net264),
    .B(\scs.oversample_in[4] ),
    .Y(_1419_));
 sky130_fd_sc_hd__o221a_1 _3422_ (.A1(_1452_),
    .A2(\scs.oversample_in[3] ),
    .B1(\scs.oversample_in[0] ),
    .B2(_1455_),
    .C1(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__o221a_1 _3423_ (.A1(net255),
    .A2(_1483_),
    .B1(_1485_),
    .B2(net270),
    .C1(_1416_),
    .X(_1421_));
 sky130_fd_sc_hd__and4_1 _3424_ (.A(_1417_),
    .B(_1418_),
    .C(_1420_),
    .D(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__and3_1 _3425_ (.A(net439),
    .B(_1415_),
    .C(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__xnor2_1 _3426_ (.A(net428),
    .B(net271),
    .Y(_1424_));
 sky130_fd_sc_hd__a211oi_1 _3427_ (.A1(_0557_),
    .A2(_1423_),
    .B1(_1424_),
    .C1(net576),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _3428_ (.A(net439),
    .B(_1454_),
    .Y(_1425_));
 sky130_fd_sc_hd__a21o_1 _3429_ (.A1(_1415_),
    .A2(_1422_),
    .B1(net240),
    .X(_1426_));
 sky130_fd_sc_hd__a21oi_1 _3430_ (.A1(net268),
    .A2(net271),
    .B1(net68),
    .Y(_1427_));
 sky130_fd_sc_hd__o221a_1 _3431_ (.A1(net268),
    .A2(net271),
    .B1(_1425_),
    .B2(_1427_),
    .C1(net513),
    .X(_0306_));
 sky130_fd_sc_hd__and3_1 _3432_ (.A(net267),
    .B(net269),
    .C(net270),
    .X(_1428_));
 sky130_fd_sc_hd__a21oi_1 _3433_ (.A1(net269),
    .A2(\scs.word_count[0] ),
    .B1(net851),
    .Y(_1429_));
 sky130_fd_sc_hd__o32a_1 _3434_ (.A1(net68),
    .A2(_1428_),
    .A3(_1429_),
    .B1(_1453_),
    .B2(net439),
    .X(_1430_));
 sky130_fd_sc_hd__nor2_1 _3435_ (.A(net581),
    .B(_1430_),
    .Y(_0307_));
 sky130_fd_sc_hd__and2_1 _3436_ (.A(net265),
    .B(_1428_),
    .X(_1431_));
 sky130_fd_sc_hd__a2bb2o_1 _3437_ (.A1_N(net67),
    .A2_N(_1431_),
    .B1(net238),
    .B2(net265),
    .X(_1432_));
 sky130_fd_sc_hd__o211a_1 _3438_ (.A1(net266),
    .A2(_1428_),
    .B1(_1432_),
    .C1(net513),
    .X(_0308_));
 sky130_fd_sc_hd__a21oi_1 _3439_ (.A1(net262),
    .A2(_1431_),
    .B1(_1426_),
    .Y(_1433_));
 sky130_fd_sc_hd__a21o_1 _3440_ (.A1(net239),
    .A2(net262),
    .B1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__o211a_1 _3441_ (.A1(net262),
    .A2(_1431_),
    .B1(_1434_),
    .C1(net511),
    .X(_0309_));
 sky130_fd_sc_hd__and3_1 _3442_ (.A(net260),
    .B(net263),
    .C(_1431_),
    .X(_1435_));
 sky130_fd_sc_hd__a2bb2o_1 _3443_ (.A1_N(net67),
    .A2_N(_1435_),
    .B1(net238),
    .B2(net261),
    .X(_1436_));
 sky130_fd_sc_hd__a31o_1 _3444_ (.A1(net262),
    .A2(net266),
    .A3(_1428_),
    .B1(net261),
    .X(_1437_));
 sky130_fd_sc_hd__and3_1 _3445_ (.A(net512),
    .B(_1436_),
    .C(_1437_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _3446_ (.A(net258),
    .B(_1435_),
    .X(_1438_));
 sky130_fd_sc_hd__a2bb2o_1 _3447_ (.A1_N(net67),
    .A2_N(_1438_),
    .B1(net238),
    .B2(net258),
    .X(_1439_));
 sky130_fd_sc_hd__o211a_1 _3448_ (.A1(net259),
    .A2(_1435_),
    .B1(_1439_),
    .C1(net512),
    .X(_0311_));
 sky130_fd_sc_hd__and3_1 _3449_ (.A(net256),
    .B(net259),
    .C(_1435_),
    .X(_1440_));
 sky130_fd_sc_hd__a2bb2o_1 _3450_ (.A1_N(net67),
    .A2_N(_1440_),
    .B1(net238),
    .B2(net256),
    .X(_1441_));
 sky130_fd_sc_hd__o211a_1 _3451_ (.A1(net257),
    .A2(_1438_),
    .B1(_1441_),
    .C1(net511),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _3452_ (.A(net255),
    .B(_1440_),
    .X(_1442_));
 sky130_fd_sc_hd__nor2_1 _3453_ (.A(net255),
    .B(_1440_),
    .Y(_1443_));
 sky130_fd_sc_hd__o32a_1 _3454_ (.A1(net68),
    .A2(_1442_),
    .A3(_1443_),
    .B1(_1449_),
    .B2(net439),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _3455_ (.A(net577),
    .B(_1444_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21oi_1 _3456_ (.A1(net427),
    .A2(_1442_),
    .B1(net254),
    .Y(_1445_));
 sky130_fd_sc_hd__a311o_1 _3457_ (.A1(net254),
    .A2(net427),
    .A3(_1442_),
    .B1(_1423_),
    .C1(net577),
    .X(_1446_));
 sky130_fd_sc_hd__nor2_1 _3458_ (.A(_1445_),
    .B(_1446_),
    .Y(_0314_));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(clknet_leaf_0_clk),
    .D(_0000_),
    .Q(\startup_cnt_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(clknet_leaf_0_clk),
    .D(_0001_),
    .Q(\startup_cnt_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(clknet_leaf_0_clk),
    .D(_0002_),
    .Q(\startup_cnt_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(clknet_leaf_0_clk),
    .D(_0003_),
    .Q(\scs.data_valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(clknet_leaf_0_clk),
    .D(_0004_),
    .Q(output_en_reg));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(clknet_leaf_0_clk),
    .D(_0005_),
    .Q(\scs.oversample_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(clknet_leaf_0_clk),
    .D(_0006_),
    .Q(\scs.oversample_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(clknet_leaf_1_clk),
    .D(_0007_),
    .Q(\scs.oversample_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(clknet_leaf_2_clk),
    .D(_0008_),
    .Q(\scs.oversample_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(clknet_leaf_11_clk),
    .D(_0009_),
    .Q(\scs.oversample_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.CLK(clknet_leaf_11_clk),
    .D(_0010_),
    .Q(\scs.oversample_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.CLK(clknet_leaf_11_clk),
    .D(_0011_),
    .Q(\scs.oversample_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.CLK(clknet_leaf_11_clk),
    .D(_0012_),
    .Q(\scs.oversample_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(clknet_leaf_11_clk),
    .D(_0013_),
    .Q(\scs.oversample_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(clknet_leaf_11_clk),
    .D(_0014_),
    .Q(\scs.oversample_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(clknet_leaf_13_clk),
    .D(net13),
    .Q(\pr.genblk1[10].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(clknet_leaf_13_clk),
    .D(net613),
    .Q(\pr.genblk1[10].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(clknet_leaf_14_clk),
    .D(net22),
    .Q(\pr.genblk1[9].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(clknet_leaf_14_clk),
    .D(net615),
    .Q(\pr.genblk1[9].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(clknet_leaf_15_clk),
    .D(net21),
    .Q(\pr.genblk1[8].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(clknet_leaf_15_clk),
    .D(net620),
    .Q(\pr.genblk1[8].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(clknet_leaf_13_clk),
    .D(net20),
    .Q(\pr.genblk1[7].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(clknet_leaf_13_clk),
    .D(net617),
    .Q(\pr.genblk1[7].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(clknet_leaf_14_clk),
    .D(net19),
    .Q(\pr.genblk1[6].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(clknet_leaf_13_clk),
    .D(net619),
    .Q(\pr.genblk1[6].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(clknet_leaf_13_clk),
    .D(net18),
    .Q(\pr.genblk1[5].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(clknet_leaf_13_clk),
    .D(net616),
    .Q(\pr.genblk1[5].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(clknet_leaf_13_clk),
    .D(net17),
    .Q(\pr.genblk1[4].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(clknet_leaf_13_clk),
    .D(net611),
    .Q(\pr.genblk1[4].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(clknet_leaf_12_clk),
    .D(net16),
    .Q(\pr.genblk1[3].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(clknet_leaf_12_clk),
    .D(net610),
    .Q(\pr.genblk1[3].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(clknet_leaf_12_clk),
    .D(net15),
    .Q(\pr.genblk1[2].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(clknet_leaf_12_clk),
    .D(net618),
    .Q(\pr.genblk1[2].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(clknet_leaf_12_clk),
    .D(net14),
    .Q(\pr.genblk1[1].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(clknet_leaf_12_clk),
    .D(net614),
    .Q(\pr.genblk1[1].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(clknet_leaf_12_clk),
    .D(net12),
    .Q(\pr.genblk1[0].pd.ff_reg_0 ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(clknet_leaf_12_clk),
    .D(net612),
    .Q(\pr.genblk1[0].pd.ff_reg_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(clknet_leaf_0_clk),
    .D(_0015_),
    .Q(\scs.enable_in ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(clknet_leaf_55_clk),
    .D(_0016_),
    .Q(\scs.diff2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(clknet_leaf_55_clk),
    .D(_0017_),
    .Q(\scs.diff2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(clknet_leaf_52_clk),
    .D(_0018_),
    .Q(\scs.diff2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(clknet_leaf_54_clk),
    .D(_0019_),
    .Q(\scs.diff2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(clknet_leaf_52_clk),
    .D(_0020_),
    .Q(\scs.diff2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(clknet_leaf_52_clk),
    .D(_0021_),
    .Q(\scs.diff2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(clknet_leaf_52_clk),
    .D(_0022_),
    .Q(\scs.diff2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(clknet_leaf_52_clk),
    .D(_0023_),
    .Q(\scs.diff2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(clknet_leaf_49_clk),
    .D(_0024_),
    .Q(\scs.diff2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(clknet_leaf_49_clk),
    .D(_0025_),
    .Q(\scs.diff2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(clknet_leaf_50_clk),
    .D(_0026_),
    .Q(\scs.diff2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(clknet_leaf_48_clk),
    .D(_0027_),
    .Q(\scs.diff2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(clknet_leaf_47_clk),
    .D(_0028_),
    .Q(\scs.diff2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(clknet_leaf_47_clk),
    .D(_0029_),
    .Q(\scs.diff2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(clknet_leaf_38_clk),
    .D(_0030_),
    .Q(\scs.diff2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(clknet_leaf_47_clk),
    .D(_0031_),
    .Q(\scs.diff2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(clknet_leaf_38_clk),
    .D(_0032_),
    .Q(\scs.diff2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(clknet_leaf_38_clk),
    .D(_0033_),
    .Q(\scs.diff2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(clknet_leaf_37_clk),
    .D(_0034_),
    .Q(\scs.diff2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(clknet_leaf_37_clk),
    .D(_0035_),
    .Q(\scs.diff2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(clknet_leaf_35_clk),
    .D(_0036_),
    .Q(\scs.diff2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(clknet_leaf_35_clk),
    .D(_0037_),
    .Q(\scs.diff2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(clknet_leaf_33_clk),
    .D(_0038_),
    .Q(\scs.diff2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(clknet_leaf_35_clk),
    .D(_0039_),
    .Q(\scs.diff2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(clknet_leaf_33_clk),
    .D(_0040_),
    .Q(\scs.diff2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(clknet_leaf_33_clk),
    .D(_0041_),
    .Q(\scs.diff2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(clknet_leaf_32_clk),
    .D(_0042_),
    .Q(\scs.diff2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(clknet_leaf_30_clk),
    .D(_0043_),
    .Q(\scs.diff2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(clknet_leaf_30_clk),
    .D(_0044_),
    .Q(\scs.diff2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(clknet_leaf_30_clk),
    .D(_0045_),
    .Q(\scs.diff2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(clknet_leaf_30_clk),
    .D(_0046_),
    .Q(\scs.diff2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(clknet_leaf_30_clk),
    .D(_0047_),
    .Q(\scs.diff2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(clknet_leaf_55_clk),
    .D(_0048_),
    .Q(\scs.diff1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(clknet_leaf_55_clk),
    .D(_0049_),
    .Q(\scs.diff1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(clknet_leaf_56_clk),
    .D(_0050_),
    .Q(\scs.diff1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(clknet_leaf_56_clk),
    .D(_0051_),
    .Q(\scs.diff1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(clknet_leaf_56_clk),
    .D(_0052_),
    .Q(\scs.diff1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(clknet_leaf_56_clk),
    .D(_0053_),
    .Q(\scs.diff1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(clknet_leaf_51_clk),
    .D(_0054_),
    .Q(\scs.diff1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(clknet_leaf_51_clk),
    .D(_0055_),
    .Q(\scs.diff1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(clknet_leaf_50_clk),
    .D(_0056_),
    .Q(\scs.diff1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(clknet_leaf_45_clk),
    .D(_0057_),
    .Q(\scs.diff1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(clknet_leaf_45_clk),
    .D(_0058_),
    .Q(\scs.diff1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(clknet_leaf_45_clk),
    .D(_0059_),
    .Q(\scs.diff1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(clknet_leaf_45_clk),
    .D(_0060_),
    .Q(\scs.diff1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.CLK(clknet_leaf_45_clk),
    .D(_0061_),
    .Q(\scs.diff1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(clknet_leaf_46_clk),
    .D(_0062_),
    .Q(\scs.diff1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(clknet_leaf_46_clk),
    .D(_0063_),
    .Q(\scs.diff1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(clknet_leaf_39_clk),
    .D(_0064_),
    .Q(\scs.diff1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(clknet_leaf_39_clk),
    .D(_0065_),
    .Q(\scs.diff1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(clknet_leaf_39_clk),
    .D(_0066_),
    .Q(\scs.diff1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(clknet_leaf_39_clk),
    .D(_0067_),
    .Q(\scs.diff1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(clknet_leaf_40_clk),
    .D(_0068_),
    .Q(\scs.diff1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(clknet_leaf_40_clk),
    .D(_0069_),
    .Q(\scs.diff1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(clknet_leaf_34_clk),
    .D(_0070_),
    .Q(\scs.diff1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(clknet_leaf_34_clk),
    .D(_0071_),
    .Q(\scs.diff1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(clknet_leaf_28_clk),
    .D(_0072_),
    .Q(\scs.diff1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(clknet_leaf_28_clk),
    .D(_0073_),
    .Q(\scs.diff1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(clknet_leaf_28_clk),
    .D(_0074_),
    .Q(\scs.diff1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(clknet_leaf_29_clk),
    .D(_0075_),
    .Q(\scs.diff1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(clknet_leaf_29_clk),
    .D(_0076_),
    .Q(\scs.diff1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(clknet_leaf_29_clk),
    .D(_0077_),
    .Q(\scs.diff1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(clknet_leaf_26_clk),
    .D(_0078_),
    .Q(\scs.diff1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(clknet_leaf_26_clk),
    .D(_0079_),
    .Q(\scs.diff1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(clknet_leaf_0_clk),
    .D(_0080_),
    .Q(\scs.acc3_d2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(clknet_leaf_56_clk),
    .D(net802),
    .Q(\scs.acc3_d2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(clknet_leaf_56_clk),
    .D(_0082_),
    .Q(\scs.acc3_d2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(clknet_leaf_56_clk),
    .D(_0083_),
    .Q(\scs.acc3_d2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(clknet_leaf_56_clk),
    .D(_0084_),
    .Q(\scs.acc3_d2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(clknet_leaf_56_clk),
    .D(_0085_),
    .Q(\scs.acc3_d2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(clknet_leaf_5_clk),
    .D(_0086_),
    .Q(\scs.acc3_d2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(clknet_leaf_5_clk),
    .D(_0087_),
    .Q(\scs.acc3_d2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(clknet_leaf_44_clk),
    .D(_0088_),
    .Q(\scs.acc3_d2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(clknet_leaf_44_clk),
    .D(net822),
    .Q(\scs.acc3_d2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(clknet_leaf_44_clk),
    .D(_0090_),
    .Q(\scs.acc3_d2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(clknet_leaf_44_clk),
    .D(_0091_),
    .Q(\scs.acc3_d2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(clknet_leaf_43_clk),
    .D(_0092_),
    .Q(\scs.acc3_d2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(clknet_leaf_43_clk),
    .D(_0093_),
    .Q(\scs.acc3_d2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(clknet_leaf_43_clk),
    .D(_0094_),
    .Q(\scs.acc3_d2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(clknet_leaf_43_clk),
    .D(_0095_),
    .Q(\scs.acc3_d2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(clknet_leaf_41_clk),
    .D(_0096_),
    .Q(\scs.acc3_d2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(clknet_leaf_41_clk),
    .D(_0097_),
    .Q(\scs.acc3_d2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(clknet_leaf_41_clk),
    .D(_0098_),
    .Q(\scs.acc3_d2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(clknet_leaf_41_clk),
    .D(_0099_),
    .Q(\scs.acc3_d2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(clknet_leaf_20_clk),
    .D(_0100_),
    .Q(\scs.acc3_d2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(clknet_leaf_40_clk),
    .D(_0101_),
    .Q(\scs.acc3_d2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(clknet_leaf_20_clk),
    .D(_0102_),
    .Q(\scs.acc3_d2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(clknet_leaf_20_clk),
    .D(_0103_),
    .Q(\scs.acc3_d2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(clknet_leaf_21_clk),
    .D(_0104_),
    .Q(\scs.acc3_d2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(clknet_leaf_21_clk),
    .D(_0105_),
    .Q(\scs.acc3_d2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(clknet_leaf_27_clk),
    .D(_0106_),
    .Q(\scs.acc3_d2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(clknet_leaf_27_clk),
    .D(_0107_),
    .Q(\scs.acc3_d2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(clknet_leaf_26_clk),
    .D(_0108_),
    .Q(\scs.acc3_d2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(clknet_leaf_26_clk),
    .D(_0109_),
    .Q(\scs.acc3_d2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.CLK(clknet_leaf_25_clk),
    .D(_0110_),
    .Q(\scs.acc3_d2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(clknet_leaf_25_clk),
    .D(net794),
    .Q(\scs.acc3_d2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(clknet_leaf_1_clk),
    .D(_0112_),
    .Q(\scs.decimation_en ));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.CLK(clknet_leaf_9_clk),
    .D(_0113_),
    .Q(\scs.acc2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.CLK(clknet_leaf_9_clk),
    .D(_0114_),
    .Q(\scs.acc2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3596_ (.CLK(clknet_leaf_9_clk),
    .D(_0115_),
    .Q(\scs.acc2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3597_ (.CLK(clknet_leaf_3_clk),
    .D(_0116_),
    .Q(\scs.acc2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(clknet_leaf_3_clk),
    .D(_0117_),
    .Q(\scs.acc2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.CLK(clknet_leaf_4_clk),
    .D(_0118_),
    .Q(\scs.acc2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(clknet_leaf_4_clk),
    .D(_0119_),
    .Q(\scs.acc2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(clknet_leaf_4_clk),
    .D(_0120_),
    .Q(\scs.acc2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(clknet_leaf_6_clk),
    .D(_0121_),
    .Q(\scs.acc2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(clknet_leaf_6_clk),
    .D(_0122_),
    .Q(\scs.acc2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(clknet_leaf_6_clk),
    .D(_0123_),
    .Q(\scs.acc2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(clknet_leaf_7_clk),
    .D(_0124_),
    .Q(\scs.acc2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(clknet_leaf_8_clk),
    .D(_0125_),
    .Q(\scs.acc2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(clknet_leaf_43_clk),
    .D(_0126_),
    .Q(\scs.acc2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(clknet_leaf_42_clk),
    .D(_0127_),
    .Q(\scs.acc2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(clknet_leaf_42_clk),
    .D(_0128_),
    .Q(\scs.acc2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(clknet_leaf_42_clk),
    .D(_0129_),
    .Q(\scs.acc2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(clknet_leaf_42_clk),
    .D(_0130_),
    .Q(\scs.acc2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.CLK(clknet_leaf_18_clk),
    .D(_0131_),
    .Q(\scs.acc2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.CLK(clknet_leaf_18_clk),
    .D(_0132_),
    .Q(\scs.acc2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(clknet_leaf_19_clk),
    .D(_0133_),
    .Q(\scs.acc2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(clknet_leaf_19_clk),
    .D(_0134_),
    .Q(\scs.acc2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(clknet_leaf_17_clk),
    .D(_0135_),
    .Q(\scs.acc2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(clknet_leaf_19_clk),
    .D(_0136_),
    .Q(\scs.acc2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(clknet_leaf_22_clk),
    .D(_0137_),
    .Q(\scs.acc2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(clknet_leaf_21_clk),
    .D(_0138_),
    .Q(\scs.acc2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(clknet_leaf_23_clk),
    .D(_0139_),
    .Q(\scs.acc2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.CLK(clknet_leaf_22_clk),
    .D(_0140_),
    .Q(\scs.acc2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.CLK(clknet_leaf_23_clk),
    .D(_0141_),
    .Q(\scs.acc2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.CLK(clknet_leaf_23_clk),
    .D(_0142_),
    .Q(\scs.acc2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(clknet_leaf_24_clk),
    .D(_0143_),
    .Q(\scs.acc2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(clknet_leaf_23_clk),
    .D(_0144_),
    .Q(\scs.acc2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.CLK(clknet_leaf_10_clk),
    .D(net877),
    .Q(\scs.acc3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.CLK(clknet_leaf_10_clk),
    .D(_0146_),
    .Q(\scs.acc3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.CLK(clknet_leaf_3_clk),
    .D(_0147_),
    .Q(\scs.acc3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(clknet_leaf_3_clk),
    .D(_0148_),
    .Q(\scs.acc3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.CLK(clknet_leaf_4_clk),
    .D(_0149_),
    .Q(\scs.acc3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(clknet_leaf_4_clk),
    .D(_0150_),
    .Q(\scs.acc3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.CLK(clknet_leaf_4_clk),
    .D(_0151_),
    .Q(\scs.acc3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(clknet_leaf_5_clk),
    .D(_0152_),
    .Q(\scs.acc3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(clknet_leaf_44_clk),
    .D(_0153_),
    .Q(\scs.acc3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(clknet_leaf_5_clk),
    .D(_0154_),
    .Q(\scs.acc3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(clknet_leaf_44_clk),
    .D(_0155_),
    .Q(\scs.acc3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(clknet_leaf_44_clk),
    .D(_0156_),
    .Q(\scs.acc3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(clknet_leaf_43_clk),
    .D(_0157_),
    .Q(\scs.acc3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(clknet_leaf_43_clk),
    .D(_0158_),
    .Q(\scs.acc3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(clknet_leaf_41_clk),
    .D(_0159_),
    .Q(\scs.acc3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(clknet_leaf_43_clk),
    .D(_0160_),
    .Q(\scs.acc3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(clknet_leaf_41_clk),
    .D(_0161_),
    .Q(\scs.acc3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(clknet_leaf_41_clk),
    .D(_0162_),
    .Q(\scs.acc3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(clknet_leaf_41_clk),
    .D(_0163_),
    .Q(\scs.acc3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(clknet_leaf_40_clk),
    .D(_0164_),
    .Q(\scs.acc3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(clknet_leaf_20_clk),
    .D(_0165_),
    .Q(\scs.acc3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(clknet_leaf_20_clk),
    .D(_0166_),
    .Q(\scs.acc3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(clknet_leaf_20_clk),
    .D(_0167_),
    .Q(\scs.acc3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(clknet_leaf_20_clk),
    .D(_0168_),
    .Q(\scs.acc3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(clknet_leaf_21_clk),
    .D(_0169_),
    .Q(\scs.acc3[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(clknet_leaf_21_clk),
    .D(_0170_),
    .Q(\scs.acc3[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_27_clk),
    .D(_0171_),
    .Q(\scs.acc3[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_21_clk),
    .D(_0172_),
    .Q(\scs.acc3[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_25_clk),
    .D(_0173_),
    .Q(\scs.acc3[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_24_clk),
    .D(_0174_),
    .Q(\scs.acc3[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_25_clk),
    .D(_0175_),
    .Q(\scs.acc3[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_24_clk),
    .D(_0176_),
    .Q(\scs.acc3[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_9_clk),
    .D(_0177_),
    .Q(\scs.acc1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3659_ (.CLK(clknet_leaf_9_clk),
    .D(_0178_),
    .Q(\scs.acc1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_9_clk),
    .D(_0179_),
    .Q(\scs.acc1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_9_clk),
    .D(_0180_),
    .Q(\scs.acc1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_3_clk),
    .D(_0181_),
    .Q(\scs.acc1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_3_clk),
    .D(net868),
    .Q(\scs.acc1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_7_clk),
    .D(_0183_),
    .Q(\scs.acc1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_7_clk),
    .D(_0184_),
    .Q(\scs.acc1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_7_clk),
    .D(_0185_),
    .Q(\scs.acc1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_7_clk),
    .D(_0186_),
    .Q(\scs.acc1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_7_clk),
    .D(_0187_),
    .Q(\scs.acc1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_8_clk),
    .D(_0188_),
    .Q(\scs.acc1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_8_clk),
    .D(_0189_),
    .Q(\scs.acc1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_8_clk),
    .D(_0190_),
    .Q(\scs.acc1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_42_clk),
    .D(_0191_),
    .Q(\scs.acc1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_42_clk),
    .D(_0192_),
    .Q(\scs.acc1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_18_clk),
    .D(_0193_),
    .Q(\scs.acc1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_18_clk),
    .D(_0194_),
    .Q(\scs.acc1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(clknet_leaf_18_clk),
    .D(_0195_),
    .Q(\scs.acc1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(clknet_leaf_18_clk),
    .D(_0196_),
    .Q(\scs.acc1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_19_clk),
    .D(_0197_),
    .Q(\scs.acc1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_17_clk),
    .D(_0198_),
    .Q(\scs.acc1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_17_clk),
    .D(_0199_),
    .Q(\scs.acc1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_16_clk),
    .D(_0200_),
    .Q(\scs.acc1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_22_clk),
    .D(_0201_),
    .Q(\scs.acc1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_22_clk),
    .D(_0202_),
    .Q(\scs.acc1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(clknet_leaf_16_clk),
    .D(_0203_),
    .Q(\scs.acc1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_22_clk),
    .D(_0204_),
    .Q(\scs.acc1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_23_clk),
    .D(_0205_),
    .Q(\scs.acc1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_23_clk),
    .D(_0206_),
    .Q(\scs.acc1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_24_clk),
    .D(_0207_),
    .Q(\scs.acc1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_16_clk),
    .D(net656),
    .Q(\scs.acc1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_54_clk),
    .D(_0209_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_54_clk),
    .D(_0210_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_53_clk),
    .D(_0211_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_54_clk),
    .D(_0212_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_53_clk),
    .D(_0213_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_53_clk),
    .D(_0214_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_53_clk),
    .D(_0215_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_53_clk),
    .D(_0216_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_49_clk),
    .D(_0217_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_48_clk),
    .D(_0218_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_48_clk),
    .D(_0219_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_48_clk),
    .D(_0220_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_48_clk),
    .D(_0221_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_47_clk),
    .D(_0222_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_47_clk),
    .D(_0223_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_38_clk),
    .D(_0224_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_38_clk),
    .D(_0225_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_38_clk),
    .D(_0226_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_37_clk),
    .D(_0227_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_37_clk),
    .D(_0228_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_36_clk),
    .D(_0229_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_36_clk),
    .D(_0230_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_36_clk),
    .D(_0231_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_36_clk),
    .D(_0232_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_33_clk),
    .D(_0233_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_32_clk),
    .D(_0234_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_32_clk),
    .D(_0235_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_32_clk),
    .D(_0236_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_31_clk),
    .D(_0237_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_31_clk),
    .D(_0238_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_31_clk),
    .D(_0239_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_31_clk),
    .D(_0240_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_55_clk),
    .D(_0241_),
    .Q(\scs.diff1_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_55_clk),
    .D(net694),
    .Q(\scs.diff1_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_55_clk),
    .D(net669),
    .Q(\scs.diff1_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_55_clk),
    .D(net679),
    .Q(\scs.diff1_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_56_clk),
    .D(net703),
    .Q(\scs.diff1_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_51_clk),
    .D(net743),
    .Q(\scs.diff1_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_51_clk),
    .D(net705),
    .Q(\scs.diff1_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_51_clk),
    .D(_0248_),
    .Q(\scs.diff1_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_50_clk),
    .D(net677),
    .Q(\scs.diff1_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_50_clk),
    .D(net671),
    .Q(\scs.diff1_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_45_clk),
    .D(_0251_),
    .Q(\scs.diff1_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_45_clk),
    .D(_0252_),
    .Q(\scs.diff1_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_46_clk),
    .D(net717),
    .Q(\scs.diff1_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_46_clk),
    .D(net773),
    .Q(\scs.diff1_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_46_clk),
    .D(net732),
    .Q(\scs.diff1_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_46_clk),
    .D(_0256_),
    .Q(\scs.diff1_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_39_clk),
    .D(net683),
    .Q(\scs.diff1_d[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_39_clk),
    .D(_0258_),
    .Q(\scs.diff1_d[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_39_clk),
    .D(_0259_),
    .Q(\scs.diff1_d[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_39_clk),
    .D(_0260_),
    .Q(\scs.diff1_d[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_39_clk),
    .D(net666),
    .Q(\scs.diff1_d[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_34_clk),
    .D(net818),
    .Q(\scs.diff1_d[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_34_clk),
    .D(net754),
    .Q(\scs.diff1_d[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_34_clk),
    .D(_0264_),
    .Q(\scs.diff1_d[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_34_clk),
    .D(net687),
    .Q(\scs.diff1_d[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_34_clk),
    .D(net689),
    .Q(\scs.diff1_d[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_28_clk),
    .D(net836),
    .Q(\scs.diff1_d[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_28_clk),
    .D(net849),
    .Q(\scs.diff1_d[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_29_clk),
    .D(net766),
    .Q(\scs.diff1_d[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_29_clk),
    .D(net727),
    .Q(\scs.diff1_d[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_29_clk),
    .D(net721),
    .Q(\scs.diff1_d[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_29_clk),
    .D(net662),
    .Q(\scs.diff1_d[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_54_clk),
    .D(_0273_),
    .Q(\scs.diff2_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_55_clk),
    .D(net700),
    .Q(\scs.diff2_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_54_clk),
    .D(net736),
    .Q(\scs.diff2_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_54_clk),
    .D(net757),
    .Q(\scs.diff2_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_53_clk),
    .D(net673),
    .Q(\scs.diff2_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_53_clk),
    .D(net723),
    .Q(\scs.diff2_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_52_clk),
    .D(net698),
    .Q(\scs.diff2_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_53_clk),
    .D(net829),
    .Q(\scs.diff2_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_49_clk),
    .D(net681),
    .Q(\scs.diff2_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_49_clk),
    .D(net729),
    .Q(\scs.diff2_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_48_clk),
    .D(net692),
    .Q(\scs.diff2_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_48_clk),
    .D(net675),
    .Q(\scs.diff2_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_47_clk),
    .D(_0285_),
    .Q(\scs.diff2_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_47_clk),
    .D(net764),
    .Q(\scs.diff2_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_47_clk),
    .D(net622),
    .Q(\scs.diff2_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_47_clk),
    .D(_0288_),
    .Q(\scs.diff2_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_38_clk),
    .D(net725),
    .Q(\scs.diff2_d[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_38_clk),
    .D(_0290_),
    .Q(\scs.diff2_d[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(clknet_leaf_37_clk),
    .D(_0291_),
    .Q(\scs.diff2_d[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(clknet_leaf_37_clk),
    .D(_0292_),
    .Q(\scs.diff2_d[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(clknet_leaf_35_clk),
    .D(net719),
    .Q(\scs.diff2_d[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(clknet_leaf_35_clk),
    .D(_0294_),
    .Q(\scs.diff2_d[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(clknet_leaf_35_clk),
    .D(net786),
    .Q(\scs.diff2_d[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(clknet_leaf_33_clk),
    .D(net685),
    .Q(\scs.diff2_d[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(clknet_leaf_33_clk),
    .D(_0297_),
    .Q(\scs.diff2_d[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(clknet_leaf_33_clk),
    .D(net714),
    .Q(\scs.diff2_d[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(clknet_leaf_32_clk),
    .D(net832),
    .Q(\scs.diff2_d[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(clknet_leaf_32_clk),
    .D(net847),
    .Q(\scs.diff2_d[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(clknet_leaf_30_clk),
    .D(net745),
    .Q(\scs.diff2_d[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(clknet_leaf_31_clk),
    .D(net784),
    .Q(\scs.diff2_d[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(clknet_leaf_30_clk),
    .D(net778),
    .Q(\scs.diff2_d[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(clknet_leaf_30_clk),
    .D(net708),
    .Q(\scs.diff2_d[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(clknet_leaf_1_clk),
    .D(_0305_),
    .Q(\scs.word_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(clknet_leaf_2_clk),
    .D(_0306_),
    .Q(\scs.word_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(clknet_leaf_2_clk),
    .D(_0307_),
    .Q(\scs.word_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(clknet_leaf_10_clk),
    .D(_0308_),
    .Q(\scs.word_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(clknet_leaf_10_clk),
    .D(_0309_),
    .Q(\scs.word_count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(clknet_leaf_10_clk),
    .D(_0310_),
    .Q(\scs.word_count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(clknet_leaf_11_clk),
    .D(_0311_),
    .Q(\scs.word_count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(clknet_leaf_11_clk),
    .D(_0312_),
    .Q(\scs.word_count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(clknet_leaf_1_clk),
    .D(_0313_),
    .Q(\scs.word_count[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(clknet_leaf_1_clk),
    .D(_0314_),
    .Q(\scs.word_count[9] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_1 fanout1 (.A(\scs.acc3[30] ),
    .X(net695));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout100 (.A(net105),
    .X(net100));
 sky130_fd_sc_hd__buf_1 fanout101 (.A(net105),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_1 fanout103 (.A(net105),
    .X(net103));
 sky130_fd_sc_hd__buf_1 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_1 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_1 fanout107 (.A(net148),
    .X(net107));
 sky130_fd_sc_hd__buf_1 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout109 (.A(net111),
    .X(net109));
 sky130_fd_sc_hd__buf_1 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout111 (.A(net114),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__buf_1 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_1 fanout114 (.A(net122),
    .X(net114));
 sky130_fd_sc_hd__buf_1 fanout115 (.A(net118),
    .X(net115));
 sky130_fd_sc_hd__buf_1 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__buf_1 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_1 fanout118 (.A(net121),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net121),
    .X(net119));
 sky130_fd_sc_hd__buf_1 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_1 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_1 fanout122 (.A(net147),
    .X(net122));
 sky130_fd_sc_hd__buf_1 fanout123 (.A(net125),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout125 (.A(net133),
    .X(net125));
 sky130_fd_sc_hd__buf_1 fanout126 (.A(net133),
    .X(net126));
 sky130_fd_sc_hd__buf_1 fanout127 (.A(net130),
    .X(net127));
 sky130_fd_sc_hd__buf_1 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net132),
    .X(net129));
 sky130_fd_sc_hd__buf_1 fanout130 (.A(net132),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_1 fanout133 (.A(net146),
    .X(net133));
 sky130_fd_sc_hd__buf_1 fanout134 (.A(net136),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout136 (.A(net145),
    .X(net136));
 sky130_fd_sc_hd__buf_1 fanout137 (.A(net145),
    .X(net137));
 sky130_fd_sc_hd__buf_1 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__buf_1 fanout139 (.A(net144),
    .X(net139));
 sky130_fd_sc_hd__buf_1 fanout140 (.A(net144),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout141 (.A(net144),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_1 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_1 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_1 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_1 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout148 (.A(_1497_),
    .X(net148));
 sky130_fd_sc_hd__buf_1 fanout149 (.A(net152),
    .X(net149));
 sky130_fd_sc_hd__buf_1 fanout150 (.A(net152),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_1 fanout152 (.A(net155),
    .X(net152));
 sky130_fd_sc_hd__buf_1 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_1 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_1 fanout155 (.A(net160),
    .X(net155));
 sky130_fd_sc_hd__buf_1 fanout156 (.A(net159),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__buf_1 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_1 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_1 fanout160 (.A(net170),
    .X(net160));
 sky130_fd_sc_hd__buf_1 fanout161 (.A(net165),
    .X(net161));
 sky130_fd_sc_hd__buf_1 fanout162 (.A(net165),
    .X(net162));
 sky130_fd_sc_hd__buf_1 fanout163 (.A(net165),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_1 fanout165 (.A(net169),
    .X(net165));
 sky130_fd_sc_hd__buf_1 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__buf_1 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_1 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_1 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_1 fanout170 (.A(net192),
    .X(net170));
 sky130_fd_sc_hd__buf_1 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_1 fanout172 (.A(net175),
    .X(net172));
 sky130_fd_sc_hd__buf_1 fanout173 (.A(net175),
    .X(net173));
 sky130_fd_sc_hd__buf_1 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout175 (.A(net181),
    .X(net175));
 sky130_fd_sc_hd__buf_1 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_1 fanout177 (.A(net180),
    .X(net177));
 sky130_fd_sc_hd__buf_1 fanout178 (.A(net180),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_1 fanout181 (.A(net191),
    .X(net181));
 sky130_fd_sc_hd__buf_1 fanout182 (.A(net184),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_1 fanout184 (.A(net190),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 fanout185 (.A(net190),
    .X(net185));
 sky130_fd_sc_hd__buf_1 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__buf_1 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_1 fanout188 (.A(net190),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_1 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_1 fanout192 (.A(net235),
    .X(net192));
 sky130_fd_sc_hd__buf_1 fanout193 (.A(net196),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 fanout194 (.A(net196),
    .X(net194));
 sky130_fd_sc_hd__buf_1 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout196 (.A(net202),
    .X(net196));
 sky130_fd_sc_hd__buf_1 fanout197 (.A(net201),
    .X(net197));
 sky130_fd_sc_hd__buf_1 fanout198 (.A(net201),
    .X(net198));
 sky130_fd_sc_hd__buf_1 fanout199 (.A(net201),
    .X(net199));
 sky130_fd_sc_hd__buf_1 fanout2 (.A(\startup_cnt_reg[0] ),
    .X(net805));
 sky130_fd_sc_hd__buf_1 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_1 fanout202 (.A(net212),
    .X(net202));
 sky130_fd_sc_hd__buf_1 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__buf_1 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_1 fanout205 (.A(net211),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 fanout206 (.A(net211),
    .X(net206));
 sky130_fd_sc_hd__buf_1 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_1 fanout208 (.A(net210),
    .X(net208));
 sky130_fd_sc_hd__buf_1 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_1 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_1 fanout212 (.A(net234),
    .X(net212));
 sky130_fd_sc_hd__buf_1 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_1 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_1 fanout215 (.A(net222),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 fanout216 (.A(net222),
    .X(net216));
 sky130_fd_sc_hd__buf_1 fanout217 (.A(net221),
    .X(net217));
 sky130_fd_sc_hd__buf_1 fanout218 (.A(net221),
    .X(net218));
 sky130_fd_sc_hd__buf_1 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__buf_1 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_1 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_1 fanout222 (.A(net233),
    .X(net222));
 sky130_fd_sc_hd__buf_1 fanout223 (.A(net225),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_1 fanout225 (.A(net232),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 fanout226 (.A(net232),
    .X(net226));
 sky130_fd_sc_hd__buf_1 fanout227 (.A(net231),
    .X(net227));
 sky130_fd_sc_hd__buf_1 fanout228 (.A(net231),
    .X(net228));
 sky130_fd_sc_hd__buf_1 fanout229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__buf_1 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_1 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_1 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_1 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 fanout235 (.A(_1496_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net242),
    .X(net236));
 sky130_fd_sc_hd__buf_1 fanout237 (.A(net242),
    .X(net237));
 sky130_fd_sc_hd__buf_1 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_1 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_1 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_1 fanout242 (.A(net246),
    .X(net242));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout243 (.A(net245),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_1 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_1 fanout246 (.A(net253),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(net252),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_1 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(_1448_),
    .X(net253));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout254 (.A(\scs.word_count[9] ),
    .X(net254));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout255 (.A(\scs.word_count[8] ),
    .X(net255));
 sky130_fd_sc_hd__buf_1 fanout256 (.A(\scs.word_count[7] ),
    .X(net256));
 sky130_fd_sc_hd__buf_1 fanout257 (.A(net874),
    .X(net257));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout258 (.A(\scs.word_count[6] ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 fanout259 (.A(net837),
    .X(net259));
 sky130_fd_sc_hd__buf_1 fanout260 (.A(\scs.word_count[5] ),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 fanout261 (.A(\scs.word_count[5] ),
    .X(net261));
 sky130_fd_sc_hd__buf_1 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout264 (.A(\scs.word_count[4] ),
    .X(net264));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout265 (.A(\scs.word_count[3] ),
    .X(net265));
 sky130_fd_sc_hd__buf_1 fanout266 (.A(net843),
    .X(net266));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout267 (.A(\scs.word_count[2] ),
    .X(net267));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout268 (.A(\scs.word_count[1] ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 fanout269 (.A(\scs.word_count[1] ),
    .X(net269));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout271 (.A(\scs.word_count[0] ),
    .X(net271));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout272 (.A(\scs.acc1[30] ),
    .X(net272));
 sky130_fd_sc_hd__buf_1 fanout273 (.A(\scs.acc1[28] ),
    .X(net273));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout274 (.A(\scs.acc1[25] ),
    .X(net274));
 sky130_fd_sc_hd__buf_1 fanout275 (.A(\scs.acc1[24] ),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(\scs.acc1[23] ),
    .X(net276));
 sky130_fd_sc_hd__buf_1 fanout277 (.A(\scs.acc1[23] ),
    .X(net277));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout278 (.A(\scs.acc1[22] ),
    .X(net278));
 sky130_fd_sc_hd__buf_1 fanout279 (.A(net865),
    .X(net279));
 sky130_fd_sc_hd__buf_1 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_1 fanout281 (.A(\scs.acc1[18] ),
    .X(net281));
 sky130_fd_sc_hd__buf_1 fanout282 (.A(\scs.acc1[16] ),
    .X(net282));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout283 (.A(\scs.acc1[15] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 fanout284 (.A(\scs.acc1[15] ),
    .X(net284));
 sky130_fd_sc_hd__buf_1 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_1 fanout287 (.A(\scs.acc1[14] ),
    .X(net287));
 sky130_fd_sc_hd__buf_1 fanout288 (.A(net290),
    .X(net288));
 sky130_fd_sc_hd__buf_1 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(\scs.acc1[13] ),
    .X(net290));
 sky130_fd_sc_hd__buf_1 fanout291 (.A(\scs.acc1[12] ),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 fanout292 (.A(net826),
    .X(net292));
 sky130_fd_sc_hd__buf_1 fanout293 (.A(\scs.acc1[10] ),
    .X(net293));
 sky130_fd_sc_hd__buf_1 fanout294 (.A(\scs.acc1[9] ),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 fanout295 (.A(\scs.acc1[9] ),
    .X(net295));
 sky130_fd_sc_hd__buf_1 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__buf_1 fanout297 (.A(\scs.acc1[8] ),
    .X(net297));
 sky130_fd_sc_hd__buf_1 fanout298 (.A(\scs.acc1[6] ),
    .X(net298));
 sky130_fd_sc_hd__buf_1 fanout299 (.A(net842),
    .X(net299));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout300 (.A(\scs.acc1[5] ),
    .X(net300));
 sky130_fd_sc_hd__buf_1 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_1 fanout303 (.A(\scs.acc1[4] ),
    .X(net303));
 sky130_fd_sc_hd__buf_1 fanout304 (.A(\scs.acc1[3] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 fanout305 (.A(\scs.acc1[3] ),
    .X(net305));
 sky130_fd_sc_hd__buf_1 fanout306 (.A(\scs.acc1[2] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 fanout307 (.A(\scs.acc1[2] ),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(\scs.acc1[1] ),
    .X(net308));
 sky130_fd_sc_hd__buf_1 fanout309 (.A(\scs.acc3[29] ),
    .X(net309));
 sky130_fd_sc_hd__buf_1 fanout310 (.A(\scs.acc3[28] ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(\scs.acc3[27] ),
    .X(net311));
 sky130_fd_sc_hd__buf_1 fanout312 (.A(\scs.acc3[27] ),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 fanout313 (.A(\scs.acc3[26] ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 fanout314 (.A(\scs.acc3[26] ),
    .X(net314));
 sky130_fd_sc_hd__buf_1 fanout315 (.A(\scs.acc3[25] ),
    .X(net315));
 sky130_fd_sc_hd__buf_1 fanout316 (.A(\scs.acc3[24] ),
    .X(net316));
 sky130_fd_sc_hd__buf_1 fanout317 (.A(\scs.acc3[24] ),
    .X(net317));
 sky130_fd_sc_hd__buf_1 fanout318 (.A(\scs.acc3[23] ),
    .X(net318));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout319 (.A(net807),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 fanout320 (.A(\scs.acc3[22] ),
    .X(net320));
 sky130_fd_sc_hd__buf_1 fanout321 (.A(\scs.acc3[21] ),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 fanout322 (.A(\scs.acc3[21] ),
    .X(net322));
 sky130_fd_sc_hd__buf_1 fanout323 (.A(\scs.acc3[20] ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 fanout324 (.A(\scs.acc3[20] ),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(\scs.acc3[19] ),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 fanout326 (.A(\scs.acc3[19] ),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 fanout327 (.A(\scs.acc3[18] ),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 fanout328 (.A(\scs.acc3[18] ),
    .X(net328));
 sky130_fd_sc_hd__buf_1 fanout329 (.A(\scs.acc3[17] ),
    .X(net329));
 sky130_fd_sc_hd__buf_1 fanout330 (.A(\scs.acc3[17] ),
    .X(net330));
 sky130_fd_sc_hd__buf_1 fanout331 (.A(\scs.acc3[16] ),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 fanout332 (.A(\scs.acc3[16] ),
    .X(net332));
 sky130_fd_sc_hd__buf_2 fanout333 (.A(\scs.acc3[15] ),
    .X(net333));
 sky130_fd_sc_hd__buf_1 fanout334 (.A(\scs.acc3[15] ),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(\scs.acc3[14] ),
    .X(net335));
 sky130_fd_sc_hd__buf_1 fanout336 (.A(\scs.acc3[14] ),
    .X(net336));
 sky130_fd_sc_hd__buf_1 fanout337 (.A(\scs.acc3[13] ),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 fanout338 (.A(\scs.acc3[13] ),
    .X(net338));
 sky130_fd_sc_hd__buf_1 fanout339 (.A(\scs.acc3[12] ),
    .X(net339));
 sky130_fd_sc_hd__buf_1 fanout340 (.A(\scs.acc3[12] ),
    .X(net340));
 sky130_fd_sc_hd__buf_1 fanout341 (.A(\scs.acc3[11] ),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 fanout342 (.A(\scs.acc3[11] ),
    .X(net342));
 sky130_fd_sc_hd__buf_1 fanout343 (.A(\scs.acc3[10] ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 fanout344 (.A(net839),
    .X(net344));
 sky130_fd_sc_hd__buf_1 fanout345 (.A(\scs.acc3[9] ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 fanout346 (.A(\scs.acc3[9] ),
    .X(net346));
 sky130_fd_sc_hd__buf_1 fanout347 (.A(\scs.acc3[8] ),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 fanout348 (.A(\scs.acc3[8] ),
    .X(net348));
 sky130_fd_sc_hd__buf_1 fanout349 (.A(\scs.acc3[7] ),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 fanout350 (.A(\scs.acc3[7] ),
    .X(net350));
 sky130_fd_sc_hd__buf_1 fanout351 (.A(\scs.acc3[6] ),
    .X(net351));
 sky130_fd_sc_hd__buf_1 fanout352 (.A(\scs.acc3[6] ),
    .X(net352));
 sky130_fd_sc_hd__buf_1 fanout353 (.A(\scs.acc3[5] ),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 fanout354 (.A(\scs.acc3[5] ),
    .X(net354));
 sky130_fd_sc_hd__buf_1 fanout355 (.A(\scs.acc3[4] ),
    .X(net355));
 sky130_fd_sc_hd__buf_1 fanout356 (.A(\scs.acc3[4] ),
    .X(net356));
 sky130_fd_sc_hd__buf_1 fanout357 (.A(\scs.acc3[3] ),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 fanout358 (.A(\scs.acc3[2] ),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(\scs.acc3[1] ),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 fanout360 (.A(net816),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 fanout361 (.A(\scs.acc3[0] ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 fanout362 (.A(\scs.acc3[0] ),
    .X(net362));
 sky130_fd_sc_hd__buf_1 fanout363 (.A(\scs.acc2[30] ),
    .X(net363));
 sky130_fd_sc_hd__buf_1 fanout364 (.A(\scs.acc2[29] ),
    .X(net364));
 sky130_fd_sc_hd__buf_1 fanout365 (.A(\scs.acc2[28] ),
    .X(net365));
 sky130_fd_sc_hd__buf_1 fanout366 (.A(\scs.acc2[27] ),
    .X(net366));
 sky130_fd_sc_hd__buf_1 fanout367 (.A(\scs.acc2[27] ),
    .X(net367));
 sky130_fd_sc_hd__buf_1 fanout368 (.A(\scs.acc2[26] ),
    .X(net368));
 sky130_fd_sc_hd__buf_1 fanout369 (.A(\scs.acc2[25] ),
    .X(net369));
 sky130_fd_sc_hd__buf_1 fanout370 (.A(net856),
    .X(net370));
 sky130_fd_sc_hd__buf_1 fanout371 (.A(\scs.acc2[24] ),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 fanout372 (.A(net873),
    .X(net372));
 sky130_fd_sc_hd__buf_1 fanout373 (.A(\scs.acc2[23] ),
    .X(net373));
 sky130_fd_sc_hd__buf_1 fanout374 (.A(net878),
    .X(net374));
 sky130_fd_sc_hd__buf_1 fanout375 (.A(\scs.acc2[22] ),
    .X(net375));
 sky130_fd_sc_hd__buf_1 fanout376 (.A(net838),
    .X(net376));
 sky130_fd_sc_hd__buf_1 fanout377 (.A(\scs.acc2[21] ),
    .X(net377));
 sky130_fd_sc_hd__buf_1 fanout378 (.A(\scs.acc2[20] ),
    .X(net378));
 sky130_fd_sc_hd__buf_1 fanout379 (.A(\scs.acc2[19] ),
    .X(net379));
 sky130_fd_sc_hd__buf_1 fanout380 (.A(net879),
    .X(net380));
 sky130_fd_sc_hd__buf_1 fanout381 (.A(\scs.acc2[18] ),
    .X(net381));
 sky130_fd_sc_hd__buf_1 fanout382 (.A(\scs.acc2[17] ),
    .X(net382));
 sky130_fd_sc_hd__buf_1 fanout383 (.A(\scs.acc2[17] ),
    .X(net383));
 sky130_fd_sc_hd__buf_1 fanout384 (.A(\scs.acc2[16] ),
    .X(net384));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout385 (.A(\scs.acc2[15] ),
    .X(net385));
 sky130_fd_sc_hd__buf_1 fanout386 (.A(\scs.acc2[15] ),
    .X(net386));
 sky130_fd_sc_hd__buf_1 fanout387 (.A(\scs.acc2[14] ),
    .X(net387));
 sky130_fd_sc_hd__buf_1 fanout388 (.A(\scs.acc2[14] ),
    .X(net388));
 sky130_fd_sc_hd__buf_1 fanout389 (.A(\scs.acc2[13] ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 fanout390 (.A(\scs.acc2[13] ),
    .X(net390));
 sky130_fd_sc_hd__buf_1 fanout391 (.A(\scs.acc2[12] ),
    .X(net391));
 sky130_fd_sc_hd__buf_1 fanout392 (.A(\scs.acc2[12] ),
    .X(net392));
 sky130_fd_sc_hd__buf_1 fanout393 (.A(\scs.acc2[11] ),
    .X(net393));
 sky130_fd_sc_hd__buf_1 fanout394 (.A(\scs.acc2[10] ),
    .X(net394));
 sky130_fd_sc_hd__buf_1 fanout395 (.A(\scs.acc2[9] ),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 fanout396 (.A(\scs.acc2[9] ),
    .X(net396));
 sky130_fd_sc_hd__buf_1 fanout397 (.A(\scs.acc2[8] ),
    .X(net397));
 sky130_fd_sc_hd__buf_1 fanout398 (.A(\scs.acc2[8] ),
    .X(net398));
 sky130_fd_sc_hd__buf_1 fanout399 (.A(\scs.acc2[7] ),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 fanout400 (.A(\scs.acc2[7] ),
    .X(net400));
 sky130_fd_sc_hd__buf_1 fanout401 (.A(\scs.acc2[6] ),
    .X(net401));
 sky130_fd_sc_hd__buf_1 fanout402 (.A(\scs.acc2[6] ),
    .X(net402));
 sky130_fd_sc_hd__buf_1 fanout403 (.A(\scs.acc2[5] ),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 fanout404 (.A(\scs.acc2[5] ),
    .X(net404));
 sky130_fd_sc_hd__buf_1 fanout405 (.A(\scs.acc2[4] ),
    .X(net405));
 sky130_fd_sc_hd__buf_1 fanout406 (.A(\scs.acc2[4] ),
    .X(net406));
 sky130_fd_sc_hd__buf_1 fanout407 (.A(\scs.acc2[3] ),
    .X(net407));
 sky130_fd_sc_hd__buf_1 fanout408 (.A(\scs.acc2[3] ),
    .X(net408));
 sky130_fd_sc_hd__buf_1 fanout409 (.A(\scs.acc2[2] ),
    .X(net409));
 sky130_fd_sc_hd__buf_1 fanout410 (.A(\scs.acc2[2] ),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 fanout411 (.A(\scs.acc2[1] ),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(\scs.acc2[0] ),
    .X(net412));
 sky130_fd_sc_hd__buf_1 fanout413 (.A(\scs.diff1[21] ),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 fanout414 (.A(\scs.diff1[19] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 fanout415 (.A(\scs.diff1[18] ),
    .X(net415));
 sky130_fd_sc_hd__buf_1 fanout416 (.A(\scs.diff1[17] ),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(\scs.diff1[15] ),
    .X(net417));
 sky130_fd_sc_hd__buf_1 fanout418 (.A(\scs.diff1[7] ),
    .X(net418));
 sky130_fd_sc_hd__buf_1 fanout419 (.A(\scs.diff2[21] ),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_2 fanout420 (.A(\scs.diff2[19] ),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(\scs.diff2[18] ),
    .X(net421));
 sky130_fd_sc_hd__buf_1 fanout422 (.A(\scs.diff2[17] ),
    .X(net422));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout423 (.A(\scs.diff2[15] ),
    .X(net423));
 sky130_fd_sc_hd__buf_1 fanout424 (.A(\scs.diff2[7] ),
    .X(net424));
 sky130_fd_sc_hd__buf_1 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 fanout426 (.A(net429),
    .X(net426));
 sky130_fd_sc_hd__buf_1 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_1 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_1 fanout429 (.A(net433),
    .X(net429));
 sky130_fd_sc_hd__buf_1 fanout430 (.A(net432),
    .X(net430));
 sky130_fd_sc_hd__buf_1 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_1 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_1 fanout433 (.A(net440),
    .X(net433));
 sky130_fd_sc_hd__buf_1 fanout434 (.A(net437),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 fanout435 (.A(net437),
    .X(net435));
 sky130_fd_sc_hd__buf_1 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_1 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_1 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__buf_1 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout440 (.A(net453),
    .X(net440));
 sky130_fd_sc_hd__buf_1 fanout441 (.A(net448),
    .X(net441));
 sky130_fd_sc_hd__buf_1 fanout442 (.A(net448),
    .X(net442));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout443 (.A(net447),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 fanout444 (.A(net447),
    .X(net444));
 sky130_fd_sc_hd__buf_1 fanout445 (.A(net447),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 fanout446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_1 fanout448 (.A(net452),
    .X(net448));
 sky130_fd_sc_hd__buf_1 fanout449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__buf_1 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_1 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_1 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_1 fanout453 (.A(net471),
    .X(net453));
 sky130_fd_sc_hd__buf_1 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 fanout455 (.A(net459),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 fanout456 (.A(net459),
    .X(net456));
 sky130_fd_sc_hd__buf_1 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_1 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_1 fanout459 (.A(net462),
    .X(net459));
 sky130_fd_sc_hd__buf_1 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_1 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_1 fanout462 (.A(net470),
    .X(net462));
 sky130_fd_sc_hd__buf_1 fanout463 (.A(net467),
    .X(net463));
 sky130_fd_sc_hd__buf_1 fanout464 (.A(net467),
    .X(net464));
 sky130_fd_sc_hd__buf_1 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_1 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_2 fanout467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_1 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_2 fanout471 (.A(\scs.enable_in ),
    .X(net471));
 sky130_fd_sc_hd__buf_1 fanout472 (.A(\startup_cnt_reg[1] ),
    .X(net472));
 sky130_fd_sc_hd__buf_1 fanout473 (.A(net477),
    .X(net473));
 sky130_fd_sc_hd__buf_1 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__buf_1 fanout475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__buf_1 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_1 fanout477 (.A(net482),
    .X(net477));
 sky130_fd_sc_hd__buf_1 fanout478 (.A(net480),
    .X(net478));
 sky130_fd_sc_hd__buf_1 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_1 fanout480 (.A(net482),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_1 fanout482 (.A(net490),
    .X(net482));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout484 (.A(net489),
    .X(net484));
 sky130_fd_sc_hd__buf_1 fanout485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__buf_1 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout487 (.A(net489),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_1 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_1 fanout490 (.A(net508),
    .X(net490));
 sky130_fd_sc_hd__buf_1 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_1 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_1 fanout493 (.A(net499),
    .X(net493));
 sky130_fd_sc_hd__buf_1 fanout494 (.A(net499),
    .X(net494));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout495 (.A(net497),
    .X(net495));
 sky130_fd_sc_hd__buf_1 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout497 (.A(net499),
    .X(net497));
 sky130_fd_sc_hd__buf_1 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout499 (.A(net507),
    .X(net499));
 sky130_fd_sc_hd__buf_1 fanout500 (.A(net503),
    .X(net500));
 sky130_fd_sc_hd__buf_1 fanout501 (.A(net503),
    .X(net501));
 sky130_fd_sc_hd__buf_1 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout503 (.A(net506),
    .X(net503));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout504 (.A(net506),
    .X(net504));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_1 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_1 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_1 fanout508 (.A(net521),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_2 fanout509 (.A(net515),
    .X(net509));
 sky130_fd_sc_hd__buf_1 fanout510 (.A(net515),
    .X(net510));
 sky130_fd_sc_hd__buf_1 fanout511 (.A(net513),
    .X(net511));
 sky130_fd_sc_hd__buf_1 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_1 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_2 fanout515 (.A(net520),
    .X(net515));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_2 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_2 fanout518 (.A(net520),
    .X(net518));
 sky130_fd_sc_hd__buf_1 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__buf_1 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_1 fanout521 (.A(net573),
    .X(net521));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout522 (.A(net526),
    .X(net522));
 sky130_fd_sc_hd__buf_1 fanout523 (.A(net526),
    .X(net523));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout524 (.A(net526),
    .X(net524));
 sky130_fd_sc_hd__buf_1 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout526 (.A(net529),
    .X(net526));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_1 fanout529 (.A(net535),
    .X(net529));
 sky130_fd_sc_hd__buf_1 fanout530 (.A(net534),
    .X(net530));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout531 (.A(net534),
    .X(net531));
 sky130_fd_sc_hd__buf_1 fanout532 (.A(net534),
    .X(net532));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__buf_1 fanout535 (.A(net557),
    .X(net535));
 sky130_fd_sc_hd__buf_1 fanout536 (.A(net540),
    .X(net536));
 sky130_fd_sc_hd__buf_1 fanout537 (.A(net540),
    .X(net537));
 sky130_fd_sc_hd__buf_1 fanout538 (.A(net540),
    .X(net538));
 sky130_fd_sc_hd__buf_1 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout540 (.A(net546),
    .X(net540));
 sky130_fd_sc_hd__buf_1 fanout541 (.A(net545),
    .X(net541));
 sky130_fd_sc_hd__buf_1 fanout542 (.A(net545),
    .X(net542));
 sky130_fd_sc_hd__buf_1 fanout543 (.A(net545),
    .X(net543));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__buf_1 fanout546 (.A(net556),
    .X(net546));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout547 (.A(net549),
    .X(net547));
 sky130_fd_sc_hd__buf_1 fanout548 (.A(net555),
    .X(net548));
 sky130_fd_sc_hd__buf_1 fanout549 (.A(net555),
    .X(net549));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout550 (.A(net554),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_1 fanout551 (.A(net554),
    .X(net551));
 sky130_fd_sc_hd__buf_1 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__buf_1 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_1 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__buf_1 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_1 fanout556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__buf_1 fanout557 (.A(net572),
    .X(net557));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout558 (.A(net560),
    .X(net558));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_2 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_1 fanout563 (.A(net571),
    .X(net563));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout564 (.A(net566),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout566 (.A(net569),
    .X(net566));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__buf_1 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_1 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_1 fanout57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__buf_1 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_1 fanout572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 fanout573 (.A(_1478_),
    .X(net573));
 sky130_fd_sc_hd__buf_2 fanout574 (.A(net592),
    .X(net574));
 sky130_fd_sc_hd__buf_1 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout576 (.A(net578),
    .X(net576));
 sky130_fd_sc_hd__buf_1 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_2 fanout578 (.A(net583),
    .X(net578));
 sky130_fd_sc_hd__buf_1 fanout579 (.A(net583),
    .X(net579));
 sky130_fd_sc_hd__buf_1 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_1 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout583 (.A(net591),
    .X(net583));
 sky130_fd_sc_hd__buf_1 fanout584 (.A(net587),
    .X(net584));
 sky130_fd_sc_hd__buf_1 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_2 fanout587 (.A(net590),
    .X(net587));
 sky130_fd_sc_hd__buf_1 fanout588 (.A(net590),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_1 fanout59 (.A(_1100_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_1 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(net608),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 fanout593 (.A(net607),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net598),
    .X(net594));
 sky130_fd_sc_hd__buf_1 fanout595 (.A(net598),
    .X(net595));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout596 (.A(net598),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_1 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 fanout598 (.A(net606),
    .X(net598));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_2 fanout60 (.A(_1116_),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout600 (.A(net605),
    .X(net600));
 sky130_fd_sc_hd__buf_1 fanout601 (.A(net603),
    .X(net601));
 sky130_fd_sc_hd__buf_1 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__buf_1 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_1 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_1 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_2 fanout608 (.A(net23),
    .X(net608));
 sky130_fd_sc_hd__buf_1 fanout61 (.A(_1094_),
    .X(net61));
 sky130_fd_sc_hd__buf_1 fanout62 (.A(_1094_),
    .X(net62));
 sky130_fd_sc_hd__buf_1 fanout63 (.A(_1086_),
    .X(net63));
 sky130_fd_sc_hd__buf_1 fanout64 (.A(_1239_),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout65 (.A(_0669_),
    .X(net65));
 sky130_fd_sc_hd__buf_1 fanout66 (.A(_1603_),
    .X(net66));
 sky130_fd_sc_hd__buf_1 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout68 (.A(_1426_),
    .X(net68));
 sky130_fd_sc_hd__buf_1 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_1 fanout70 (.A(_1103_),
    .X(net70));
 sky130_fd_sc_hd__buf_1 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout73 (.A(net79),
    .X(net73));
 sky130_fd_sc_hd__buf_1 fanout74 (.A(net79),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout75 (.A(net78),
    .X(net75));
 sky130_fd_sc_hd__buf_1 fanout76 (.A(net78),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_1 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_1 fanout79 (.A(net87),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout81 (.A(net86),
    .X(net81));
 sky130_fd_sc_hd__buf_1 fanout82 (.A(net85),
    .X(net82));
 sky130_fd_sc_hd__buf_1 fanout83 (.A(net85),
    .X(net83));
 sky130_fd_sc_hd__buf_1 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_1 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_1 fanout87 (.A(net107),
    .X(net87));
 sky130_fd_sc_hd__buf_1 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__buf_1 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_1 fanout91 (.A(net97),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_1 fanout93 (.A(net96),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout94 (.A(net96),
    .X(net94));
 sky130_fd_sc_hd__buf_1 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_1 fanout97 (.A(net106),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout98 (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\pr.genblk1[2].pd.ff_reg_0 ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0304_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\scs.acc3_d2[6] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\scs.diff1_d[0] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\scs.acc1[20] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\scs.acc1[7] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\scs.diff2[25] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0298_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\scs.diff1_d[11] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\scs.diff1[12] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0253_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\pr.genblk1[6].pd.ff_reg_0 ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\scs.diff2[20] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0293_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\scs.diff1[30] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0271_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\scs.diff2[5] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0278_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\scs.diff2[16] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0289_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\scs.diff1[29] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0270_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\pr.genblk1[8].pd.ff_reg_0 ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\scs.diff2[9] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0282_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\scs.diff1_d[10] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\scs.diff1[14] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0255_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\scs.diff2[12] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\scs.acc2[20] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\scs.diff2[2] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0275_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\scs.acc1[29] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\scs.diff2[14] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\scs.acc1[17] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\scs.diff2_d[12] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\scs.diff2[24] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\scs.diff2_d[24] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\scs.diff1[5] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0246_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\scs.diff2[28] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0301_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net32),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net39),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0287_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net33),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net54),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\scs.diff2[0] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\scs.diff1[0] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net42),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\scs.diff1[22] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0263_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\scs.acc3_d2[22] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\scs.diff2[3] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0276_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\scs.acc2[26] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net50),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net41),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\scs.acc3_d2[8] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\scs.acc3_d2[14] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\scs.diff2[18] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\scs.diff2[13] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0286_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\scs.diff1[28] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0269_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net29),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\scs.acc2[1] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net48),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\scs.diff2_d[0] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\scs.diff2[17] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\scs.acc3_d2[20] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\scs.diff1[13] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0254_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\scs.acc3_d2[29] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\scs.acc1[24] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\scs.acc2[16] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\scs.diff2[30] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\scs.acc2[18] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0303_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\scs.acc3_d2[25] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\scs.acc3_d2[28] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\scs.diff1[18] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\scs.acc3_d2[2] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\scs.diff2[29] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0302_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\scs.diff2[22] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0295_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\scs.acc3_d2[3] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net38),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\scs.acc3_d2[5] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\scs.acc3_d2[0] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\scs.acc3_d2[12] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\scs.acc3_d2[13] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\scs.acc3[30] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\scs.acc3_d2[31] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0111_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\scs.acc3_d2[11] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\scs.acc3_d2[30] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\scs.acc3_d2[24] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net40),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\scs.acc3_d2[23] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\scs.acc3_d2[10] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net26),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\scs.acc3_d2[1] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0081_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\scs.acc1[10] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\scs.acc3[29] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net361),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\scs.acc3[22] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\pr.genblk1[3].pd.ff_reg_0 ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net27),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\scs.diff1[17] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\scs.acc1[21] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\scs.acc3_d2[16] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\scs.acc3_d2[17] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\scs.acc3[2] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net47),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\scs.acc3[3] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\scs.diff2_d[21] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\scs.acc3[1] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\scs.diff1_d[21] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\scs.acc2[11] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0262_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\scs.acc3_d2[21] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\scs.diff1_d[17] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\scs.acc3_d2[9] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0089_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\scs.acc1[26] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\scs.diff2_d[17] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\scs.diff1_d[15] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\scs.acc1[12] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\scs.diff1_d[7] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net31),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\scs.diff2_d[7] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0280_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\scs.acc1[0] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\scs.diff2[26] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0299_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\scs.diff2_d[15] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\scs.acc3_d2[7] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\scs.diff1[26] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0267_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\scs.word_count[6] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net52),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\scs.acc2[22] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\scs.acc3[10] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\startup_cnt_reg[2] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_1486_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\scs.acc1[6] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\scs.word_count[3] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\scs.diff1_d[19] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\scs.diff2[27] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0300_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net35),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\scs.diff1_d[27] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0268_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\scs.acc3[28] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\scs.word_count[2] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net25),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\scs.diff2_d[19] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\scs.diff1[27] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\scs.acc2[25] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\startup_cnt_reg[2] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net24),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\scs.acc3_d2[15] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\scs.acc3_d2[18] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\scs.acc1[27] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\scs.acc3_d2[26] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\scs.acc3_d2[27] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\startup_cnt_reg[0] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\scs.acc3_d2[19] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\scs.acc1[19] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_1082_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net37),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0182_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net408),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net410),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\scs.acc2[24] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\scs.word_count[7] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net362),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0145_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net34),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\scs.acc2[23] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\scs.acc2[19] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0559_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\scs.decimation_en ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\scs.acc2[0] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\pr.genblk1[4].pd.ff_reg_0 ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0560_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\scs.diff2[19] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\scs.diff1[7] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net55),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net53),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net28),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net49),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net30),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net51),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net43),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\pr.genblk1[0].pd.ff_reg_0 ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net45),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net44),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\scs.diff2[21] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\scs.acc1[11] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\scs.diff1[19] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\scs.diff1[11] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\scs.diff1[21] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\scs.acc1[31] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0208_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\scs.diff2[7] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\pr.genblk1[10].pd.ff_reg_0 ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\scs.diff1[15] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\scs.diff1[23] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\scs.acc1[28] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\scs.diff1[31] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0272_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\scs.diff1_d[23] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net46),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\scs.diff1[20] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0261_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\scs.diff2[15] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\pr.genblk1[1].pd.ff_reg_0 ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\scs.diff1[2] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0243_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\scs.diff1[9] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0250_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\scs.diff2[4] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0277_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\scs.diff2[11] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0284_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\scs.diff1[8] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0249_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\pr.genblk1[9].pd.ff_reg_0 ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\scs.diff1[3] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0244_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\scs.diff2[8] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0281_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\scs.diff1[16] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0257_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\scs.diff2[23] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0296_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\scs.diff1[24] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0265_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\pr.genblk1[5].pd.ff_reg_0 ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\scs.diff1[25] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0266_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\scs.diff1[10] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\scs.diff2[10] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0283_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\scs.diff1[1] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0242_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_1712_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\scs.diff2[6] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\pr.genblk1[7].pd.ff_reg_0 ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0279_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\scs.diff2[1] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0274_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net36),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\scs.diff1[4] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0245_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\scs.diff1[6] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0247_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\scs.acc3_d2[4] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\scs.diff2[31] ),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(enable_in),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(oversample_in[8]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(oversample_in[9]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(phase_in[0]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(phase_in[10]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(phase_in[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(phase_in[2]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(phase_in[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(phase_in[4]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(phase_in[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(phase_in[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(oversample_in[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(phase_in[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(phase_in[8]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(phase_in[9]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(rst),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(oversample_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(oversample_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(oversample_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(oversample_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(oversample_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(oversample_in[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(oversample_in[7]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 output24 (.A(net24),
    .X(data_out[0]));
 sky130_fd_sc_hd__buf_1 output25 (.A(net25),
    .X(data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(data_out[11]));
 sky130_fd_sc_hd__buf_1 output27 (.A(net27),
    .X(data_out[12]));
 sky130_fd_sc_hd__buf_1 output28 (.A(net28),
    .X(data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(data_out[14]));
 sky130_fd_sc_hd__buf_1 output30 (.A(net30),
    .X(data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(data_out[16]));
 sky130_fd_sc_hd__buf_1 output32 (.A(net32),
    .X(data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(data_out[18]));
 sky130_fd_sc_hd__buf_1 output34 (.A(net34),
    .X(data_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(data_out[20]));
 sky130_fd_sc_hd__buf_1 output37 (.A(net37),
    .X(data_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(data_out[22]));
 sky130_fd_sc_hd__buf_1 output39 (.A(net39),
    .X(data_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(data_out[24]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(data_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(data_out[26]));
 sky130_fd_sc_hd__buf_1 output43 (.A(net43),
    .X(data_out[27]));
 sky130_fd_sc_hd__buf_1 output44 (.A(net44),
    .X(data_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(data_out[29]));
 sky130_fd_sc_hd__buf_1 output46 (.A(net46),
    .X(data_out[2]));
 sky130_fd_sc_hd__buf_1 output47 (.A(net47),
    .X(data_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(data_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_1 output50 (.A(net50),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_1 output52 (.A(net52),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(data_out[7]));
 sky130_fd_sc_hd__buf_1 output54 (.A(net54),
    .X(data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(data_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(data_valid_out));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(_0580_),
    .X(net609));
endmodule

