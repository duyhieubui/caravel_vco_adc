magic
tech sky130A
magscale 1 2
timestamp 1637984468
<< locali >>
rect 98653 573087 98687 573189
rect 480821 572747 480855 572917
rect 465733 401489 465917 401523
rect 465733 401455 465767 401489
rect 369133 400639 369167 401149
rect 378793 400707 378827 401421
rect 465641 400979 465675 401285
rect 177991 321589 178141 321623
rect 179705 321555 179739 321657
rect 177037 320807 177071 321317
rect 176945 320263 176979 320501
rect 177221 320399 177255 321385
rect 185593 320263 185627 320365
rect 50261 319311 50295 320025
rect 60013 319379 60047 320025
rect 177957 319719 177991 320229
rect 181085 320195 181119 320229
rect 185501 320195 185535 320229
rect 185685 320195 185719 320365
rect 181085 320161 181269 320195
rect 185501 320161 185719 320195
rect 185777 320195 185811 321521
rect 179797 320025 179889 320059
rect 179797 319311 179831 320025
rect 179889 319515 179923 319889
rect 179981 319515 180015 320093
rect 50111 319277 50295 319311
rect 179555 319277 179831 319311
rect 180073 319311 180107 319957
rect 185501 319923 185535 320025
rect 185409 319787 185443 319889
rect 185409 319753 185777 319787
rect 182005 319243 182039 319481
rect 204913 319107 204947 319753
rect 19349 286807 19383 287861
rect 19441 277355 19475 277457
rect 19993 277397 20027 286977
rect 19993 277363 20671 277397
rect 19441 258043 19475 258145
rect 19441 238731 19475 238833
rect 20637 229097 20671 277363
rect 178693 267631 178727 283033
rect 178785 282931 178819 287385
rect 180717 267737 180751 287385
rect 337853 287079 337887 288745
rect 337117 282591 337151 286841
rect 337945 286807 337979 287249
rect 179981 267703 180751 267737
rect 178693 257975 178727 258077
rect 179613 253759 179647 258009
rect 179981 257839 180015 267703
rect 179521 234719 179555 244341
rect 179981 244171 180015 253861
rect 179797 234651 179831 244001
rect 19993 229063 20671 229097
rect 19441 219419 19475 219521
rect 19441 203915 19475 209729
rect 19533 209355 19567 209661
rect 19625 209423 19659 209865
rect 19993 209831 20027 229063
rect 179429 224859 179463 225029
rect 179981 224995 180015 234685
rect 165813 203847 165847 204289
rect 165905 203779 165939 204153
rect 165997 203847 166031 204221
rect 166089 203983 166123 204221
rect 166181 204051 166215 204153
rect 175783 204085 176117 204119
rect 175657 204017 175933 204051
rect 175657 203983 175691 204017
rect 166089 203813 166457 203847
rect 166089 203779 166123 203813
rect 165905 203745 166123 203779
rect 166181 203303 166215 203473
rect 166273 203371 166307 203473
rect 178049 203099 178083 205717
rect 179613 205683 179647 215237
rect 179981 215203 180015 224825
rect 179705 203303 179739 205785
rect 181453 204017 181637 204051
rect 181453 203983 181487 204017
rect 27629 3859 27663 4029
rect 125149 2839 125183 3689
<< viali >>
rect 98653 573189 98687 573223
rect 98653 573053 98687 573087
rect 480821 572917 480855 572951
rect 480821 572713 480855 572747
rect 465917 401489 465951 401523
rect 378793 401421 378827 401455
rect 465733 401421 465767 401455
rect 369133 401149 369167 401183
rect 465641 401285 465675 401319
rect 465641 400945 465675 400979
rect 378793 400673 378827 400707
rect 369133 400605 369167 400639
rect 179705 321657 179739 321691
rect 177957 321589 177991 321623
rect 178141 321589 178175 321623
rect 179705 321521 179739 321555
rect 185777 321521 185811 321555
rect 177221 321385 177255 321419
rect 177037 321317 177071 321351
rect 177037 320773 177071 320807
rect 176945 320501 176979 320535
rect 177221 320365 177255 320399
rect 185593 320365 185627 320399
rect 176945 320229 176979 320263
rect 177957 320229 177991 320263
rect 50261 320025 50295 320059
rect 60013 320025 60047 320059
rect 181085 320229 181119 320263
rect 185501 320229 185535 320263
rect 185593 320229 185627 320263
rect 185685 320365 185719 320399
rect 181269 320161 181303 320195
rect 185777 320161 185811 320195
rect 179981 320093 180015 320127
rect 177957 319685 177991 319719
rect 179889 320025 179923 320059
rect 60013 319345 60047 319379
rect 179889 319889 179923 319923
rect 179889 319481 179923 319515
rect 185501 320025 185535 320059
rect 179981 319481 180015 319515
rect 180073 319957 180107 319991
rect 50077 319277 50111 319311
rect 179521 319277 179555 319311
rect 185409 319889 185443 319923
rect 185501 319889 185535 319923
rect 185777 319753 185811 319787
rect 204913 319753 204947 319787
rect 180073 319277 180107 319311
rect 182005 319481 182039 319515
rect 182005 319209 182039 319243
rect 204913 319073 204947 319107
rect 337853 288745 337887 288779
rect 19349 287861 19383 287895
rect 178785 287385 178819 287419
rect 19349 286773 19383 286807
rect 19993 286977 20027 287011
rect 19441 277457 19475 277491
rect 178693 283033 178727 283067
rect 19441 277321 19475 277355
rect 19441 258145 19475 258179
rect 19441 258009 19475 258043
rect 19441 238833 19475 238867
rect 19441 238697 19475 238731
rect 178785 282897 178819 282931
rect 180717 287385 180751 287419
rect 337853 287045 337887 287079
rect 337945 287249 337979 287283
rect 337117 286841 337151 286875
rect 337945 286773 337979 286807
rect 337117 282557 337151 282591
rect 178693 267597 178727 267631
rect 178693 258077 178727 258111
rect 178693 257941 178727 257975
rect 179613 258009 179647 258043
rect 179981 257805 180015 257839
rect 179613 253725 179647 253759
rect 179981 253861 180015 253895
rect 179521 244341 179555 244375
rect 179981 244137 180015 244171
rect 179521 234685 179555 234719
rect 179797 244001 179831 244035
rect 179797 234617 179831 234651
rect 179981 234685 180015 234719
rect 19441 219521 19475 219555
rect 19441 219385 19475 219419
rect 19625 209865 19659 209899
rect 19441 209729 19475 209763
rect 19533 209661 19567 209695
rect 179429 225029 179463 225063
rect 179981 224961 180015 224995
rect 179429 224825 179463 224859
rect 179981 224825 180015 224859
rect 19993 209797 20027 209831
rect 179613 215237 179647 215271
rect 19625 209389 19659 209423
rect 19533 209321 19567 209355
rect 178049 205717 178083 205751
rect 19441 203881 19475 203915
rect 165813 204289 165847 204323
rect 165997 204221 166031 204255
rect 165813 203813 165847 203847
rect 165905 204153 165939 204187
rect 166089 204221 166123 204255
rect 166181 204153 166215 204187
rect 175749 204085 175783 204119
rect 176117 204085 176151 204119
rect 166181 204017 166215 204051
rect 175933 204017 175967 204051
rect 166089 203949 166123 203983
rect 175657 203949 175691 203983
rect 165997 203813 166031 203847
rect 166457 203813 166491 203847
rect 166181 203473 166215 203507
rect 166273 203473 166307 203507
rect 166273 203337 166307 203371
rect 166181 203269 166215 203303
rect 179981 215169 180015 215203
rect 179613 205649 179647 205683
rect 179705 205785 179739 205819
rect 181637 204017 181671 204051
rect 181453 203949 181487 203983
rect 179705 203269 179739 203303
rect 178049 203065 178083 203099
rect 27629 4029 27663 4063
rect 27629 3825 27663 3859
rect 125149 3689 125183 3723
rect 125149 2805 125183 2839
<< metal1 >>
rect 332502 700952 332508 701004
rect 332560 700992 332566 701004
rect 472066 700992 472072 701004
rect 332560 700964 472072 700992
rect 332560 700952 332566 700964
rect 472066 700952 472072 700964
rect 472124 700952 472130 701004
rect 283834 700884 283840 700936
rect 283892 700924 283898 700936
rect 469214 700924 469220 700936
rect 283892 700896 469220 700924
rect 283892 700884 283898 700896
rect 469214 700884 469220 700896
rect 469272 700884 469278 700936
rect 267642 700816 267648 700868
rect 267700 700856 267706 700868
rect 470594 700856 470600 700868
rect 267700 700828 470600 700856
rect 267700 700816 267706 700828
rect 470594 700816 470600 700828
rect 470652 700816 470658 700868
rect 218974 700748 218980 700800
rect 219032 700788 219038 700800
rect 467926 700788 467932 700800
rect 219032 700760 467932 700788
rect 219032 700748 219038 700760
rect 467926 700748 467932 700760
rect 467984 700748 467990 700800
rect 202782 700680 202788 700732
rect 202840 700720 202846 700732
rect 467834 700720 467840 700732
rect 202840 700692 467840 700720
rect 202840 700680 202846 700692
rect 467834 700680 467840 700692
rect 467892 700680 467898 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 465074 700652 465080 700664
rect 154172 700624 465080 700652
rect 154172 700612 154178 700624
rect 465074 700612 465080 700624
rect 465132 700612 465138 700664
rect 56778 700544 56784 700596
rect 56836 700584 56842 700596
rect 105538 700584 105544 700596
rect 56836 700556 105544 700584
rect 56836 700544 56842 700556
rect 105538 700544 105544 700556
rect 105596 700544 105602 700596
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 466454 700584 466460 700596
rect 137888 700556 466460 700584
rect 137888 700544 137894 700556
rect 466454 700544 466460 700556
rect 466512 700544 466518 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 462222 700516 462228 700528
rect 89220 700488 462228 700516
rect 89220 700476 89226 700488
rect 462222 700476 462228 700488
rect 462280 700476 462286 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 463694 700448 463700 700460
rect 73028 700420 463700 700448
rect 73028 700408 73034 700420
rect 463694 700408 463700 700420
rect 463752 700408 463758 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 460934 700380 460940 700392
rect 24360 700352 460940 700380
rect 24360 700340 24366 700352
rect 460934 700340 460940 700352
rect 460992 700340 460998 700392
rect 462406 700380 462412 700392
rect 461688 700352 462412 700380
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 461688 700312 461716 700352
rect 462406 700340 462412 700352
rect 462464 700340 462470 700392
rect 8168 700284 461716 700312
rect 8168 700272 8174 700284
rect 462314 700272 462320 700324
rect 462372 700312 462378 700324
rect 472802 700312 472808 700324
rect 462372 700284 472808 700312
rect 462372 700272 462378 700284
rect 472802 700272 472808 700284
rect 472860 700272 472866 700324
rect 530578 700272 530584 700324
rect 530636 700312 530642 700324
rect 543458 700312 543464 700324
rect 530636 700284 543464 700312
rect 530636 700272 530642 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 348786 700204 348792 700256
rect 348844 700244 348850 700256
rect 471974 700244 471980 700256
rect 348844 700216 471980 700244
rect 348844 700204 348850 700216
rect 471974 700204 471980 700216
rect 472032 700204 472038 700256
rect 397454 700136 397460 700188
rect 397512 700176 397518 700188
rect 472710 700176 472716 700188
rect 397512 700148 472716 700176
rect 397512 700136 397518 700148
rect 472710 700136 472716 700148
rect 472768 700136 472774 700188
rect 413646 700068 413652 700120
rect 413704 700108 413710 700120
rect 472894 700108 472900 700120
rect 413704 700080 472900 700108
rect 413704 700068 413710 700080
rect 472894 700068 472900 700080
rect 472952 700068 472958 700120
rect 446122 700000 446128 700052
rect 446180 700040 446186 700052
rect 491294 700040 491300 700052
rect 446180 700012 491300 700040
rect 446180 700000 446186 700012
rect 491294 700000 491300 700012
rect 491352 700000 491358 700052
rect 250438 699660 250444 699712
rect 250496 699700 250502 699712
rect 251450 699700 251456 699712
rect 250496 699672 251456 699700
rect 250496 699660 250502 699672
rect 251450 699660 251456 699672
rect 251508 699660 251514 699712
rect 475378 699660 475384 699712
rect 475436 699700 475442 699712
rect 478506 699700 478512 699712
rect 475436 699672 478512 699700
rect 475436 699660 475442 699672
rect 478506 699660 478512 699672
rect 478564 699660 478570 699712
rect 527174 699660 527180 699712
rect 527232 699700 527238 699712
rect 528554 699700 528560 699712
rect 527232 699672 528560 699700
rect 527232 699660 527238 699672
rect 528554 699660 528560 699672
rect 528612 699660 528618 699712
rect 536098 696940 536104 696992
rect 536156 696980 536162 696992
rect 580166 696980 580172 696992
rect 536156 696952 580172 696980
rect 536156 696940 536162 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 529198 683136 529204 683188
rect 529256 683176 529262 683188
rect 580166 683176 580172 683188
rect 529256 683148 580172 683176
rect 529256 683136 529262 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 276290 682388 276296 682440
rect 276348 682428 276354 682440
rect 316034 682428 316040 682440
rect 276348 682400 316040 682428
rect 276348 682388 276354 682400
rect 316034 682388 316040 682400
rect 316092 682388 316098 682440
rect 267182 681708 267188 681760
rect 267240 681748 267246 681760
rect 276290 681748 276296 681760
rect 267240 681720 276296 681748
rect 267240 681708 267246 681720
rect 276290 681708 276296 681720
rect 276348 681748 276354 681760
rect 276750 681748 276756 681760
rect 276348 681720 276756 681748
rect 276348 681708 276354 681720
rect 276750 681708 276756 681720
rect 276808 681708 276814 681760
rect 455322 680348 455328 680400
rect 455380 680388 455386 680400
rect 483474 680388 483480 680400
rect 455380 680360 483480 680388
rect 455380 680348 455386 680360
rect 483474 680348 483480 680360
rect 483532 680348 483538 680400
rect 97902 679260 97908 679312
rect 97960 679300 97966 679312
rect 99650 679300 99656 679312
rect 97960 679272 99656 679300
rect 97960 679260 97966 679272
rect 99650 679260 99656 679272
rect 99708 679260 99714 679312
rect 241422 679260 241428 679312
rect 241480 679300 241486 679312
rect 316678 679300 316684 679312
rect 241480 679272 316684 679300
rect 241480 679260 241486 679272
rect 316678 679260 316684 679272
rect 316736 679260 316742 679312
rect 85482 678988 85488 679040
rect 85540 679028 85546 679040
rect 316770 679028 316776 679040
rect 85540 679000 316776 679028
rect 85540 678988 85546 679000
rect 316770 678988 316776 679000
rect 316828 678988 316834 679040
rect 88058 677288 88064 677340
rect 88116 677328 88122 677340
rect 93854 677328 93860 677340
rect 88116 677300 93860 677328
rect 88116 677288 88122 677300
rect 93854 677288 93860 677300
rect 93912 677288 93918 677340
rect 271874 676268 271880 676320
rect 271932 676308 271938 676320
rect 272886 676308 272892 676320
rect 271932 676280 272892 676308
rect 271932 676268 271938 676280
rect 272886 676268 272892 676280
rect 272944 676268 272950 676320
rect 78582 675452 78588 675504
rect 78640 675492 78646 675504
rect 86126 675492 86132 675504
rect 78640 675464 86132 675492
rect 78640 675452 78646 675464
rect 86126 675452 86132 675464
rect 86184 675452 86190 675504
rect 238662 675452 238668 675504
rect 238720 675492 238726 675504
rect 241514 675492 241520 675504
rect 238720 675464 241520 675492
rect 238720 675452 238726 675464
rect 241514 675452 241520 675464
rect 241572 675452 241578 675504
rect 505554 674296 505560 674348
rect 505612 674336 505618 674348
rect 506382 674336 506388 674348
rect 505612 674308 506388 674336
rect 505612 674296 505618 674308
rect 506382 674296 506388 674308
rect 506440 674296 506446 674348
rect 482922 674160 482928 674212
rect 482980 674200 482986 674212
rect 490650 674200 490656 674212
rect 482980 674172 490656 674200
rect 482980 674160 482986 674172
rect 490650 674160 490656 674172
rect 490708 674160 490714 674212
rect 477402 674092 477408 674144
rect 477460 674132 477466 674144
rect 487246 674132 487252 674144
rect 477460 674104 487252 674132
rect 477460 674092 477466 674104
rect 487246 674092 487252 674104
rect 487304 674092 487310 674144
rect 493318 673888 493324 673940
rect 493376 673928 493382 673940
rect 494422 673928 494428 673940
rect 493376 673900 494428 673928
rect 493376 673888 493382 673900
rect 494422 673888 494428 673900
rect 494480 673888 494486 673940
rect 499482 673480 499488 673532
rect 499540 673520 499546 673532
rect 500218 673520 500224 673532
rect 499540 673492 500224 673520
rect 499540 673480 499546 673492
rect 500218 673480 500224 673492
rect 500276 673480 500282 673532
rect 82722 672732 82728 672784
rect 82780 672772 82786 672784
rect 90634 672772 90640 672784
rect 82780 672744 90640 672772
rect 82780 672732 82786 672744
rect 90634 672732 90640 672744
rect 90692 672732 90698 672784
rect 92382 672732 92388 672784
rect 92440 672772 92446 672784
rect 96706 672772 96712 672784
rect 92440 672744 96712 672772
rect 92440 672732 92446 672744
rect 96706 672732 96712 672744
rect 96764 672732 96770 672784
rect 114738 672528 114744 672580
rect 114796 672568 114802 672580
rect 115842 672568 115848 672580
rect 114796 672540 115848 672568
rect 114796 672528 114802 672540
rect 115842 672528 115848 672540
rect 115900 672528 115906 672580
rect 242802 672052 242808 672104
rect 242860 672092 242866 672104
rect 246298 672092 246304 672104
rect 242860 672064 246304 672092
rect 242860 672052 242866 672064
rect 246298 672052 246304 672064
rect 246356 672052 246362 672104
rect 251174 672052 251180 672104
rect 251232 672092 251238 672104
rect 252186 672092 252192 672104
rect 251232 672064 252192 672092
rect 251232 672052 251238 672064
rect 252186 672052 252192 672064
rect 252244 672052 252250 672104
rect 258534 672052 258540 672104
rect 258592 672092 258598 672104
rect 259362 672092 259368 672104
rect 258592 672064 259368 672092
rect 258592 672052 258598 672064
rect 259362 672052 259368 672064
rect 259420 672052 259426 672104
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 323670 670732 323676 670744
rect 3568 670704 323676 670732
rect 3568 670692 3574 670704
rect 323670 670692 323676 670704
rect 323728 670692 323734 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 336090 656928 336096 656940
rect 3476 656900 336096 656928
rect 3476 656888 3482 656900
rect 336090 656888 336096 656900
rect 336148 656888 336154 656940
rect 533338 643084 533344 643136
rect 533396 643124 533402 643136
rect 580166 643124 580172 643136
rect 533396 643096 580172 643124
rect 533396 643084 533402 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 502242 632884 502248 632936
rect 502300 632924 502306 632936
rect 511442 632924 511448 632936
rect 502300 632896 511448 632924
rect 502300 632884 502306 632896
rect 511442 632884 511448 632896
rect 511500 632884 511506 632936
rect 264882 632816 264888 632868
rect 264940 632856 264946 632868
rect 272058 632856 272064 632868
rect 264940 632828 272064 632856
rect 264940 632816 264946 632828
rect 272058 632816 272064 632828
rect 272116 632816 272122 632868
rect 502426 632816 502432 632868
rect 502484 632856 502490 632868
rect 516318 632856 516324 632868
rect 502484 632828 516324 632856
rect 502484 632816 502490 632828
rect 516318 632816 516324 632828
rect 516376 632816 516382 632868
rect 270402 632748 270408 632800
rect 270460 632788 270466 632800
rect 281534 632788 281540 632800
rect 270460 632760 281540 632788
rect 270460 632748 270466 632760
rect 281534 632748 281540 632760
rect 281592 632748 281598 632800
rect 506382 632748 506388 632800
rect 506440 632788 506446 632800
rect 521286 632788 521292 632800
rect 506440 632760 521292 632788
rect 506440 632748 506446 632760
rect 521286 632748 521292 632760
rect 521344 632748 521350 632800
rect 111886 632680 111892 632732
rect 111944 632720 111950 632732
rect 116578 632720 116584 632732
rect 111944 632692 116584 632720
rect 111944 632680 111950 632692
rect 116578 632680 116584 632692
rect 116636 632680 116642 632732
rect 117682 632680 117688 632732
rect 117740 632720 117746 632732
rect 126422 632720 126428 632732
rect 117740 632692 126428 632720
rect 117740 632680 117746 632692
rect 126422 632680 126428 632692
rect 126480 632680 126486 632732
rect 271966 632680 271972 632732
rect 272024 632720 272030 632732
rect 286318 632720 286324 632732
rect 272024 632692 286324 632720
rect 272024 632680 272030 632692
rect 286318 632680 286324 632692
rect 286376 632680 286382 632732
rect 506474 632680 506480 632732
rect 506532 632720 506538 632732
rect 526162 632720 526168 632732
rect 506532 632692 526168 632720
rect 506532 632680 506538 632692
rect 526162 632680 526168 632692
rect 526220 632680 526226 632732
rect 486878 632340 486884 632392
rect 486936 632380 486942 632392
rect 491570 632380 491576 632392
rect 486936 632352 491576 632380
rect 486936 632340 486942 632352
rect 491570 632340 491576 632352
rect 491628 632340 491634 632392
rect 247678 632272 247684 632324
rect 247736 632312 247742 632324
rect 248414 632312 248420 632324
rect 247736 632284 248420 632312
rect 247736 632272 247742 632284
rect 248414 632272 248420 632284
rect 248472 632272 248478 632324
rect 260834 632136 260840 632188
rect 260892 632176 260898 632188
rect 266722 632176 266728 632188
rect 260892 632148 266728 632176
rect 260892 632136 260898 632148
rect 266722 632136 266728 632148
rect 266780 632136 266786 632188
rect 499574 632136 499580 632188
rect 499632 632176 499638 632188
rect 506566 632176 506572 632188
rect 499632 632148 506572 632176
rect 499632 632136 499638 632148
rect 506566 632136 506572 632148
rect 506624 632136 506630 632188
rect 78030 632068 78036 632120
rect 78088 632108 78094 632120
rect 78582 632108 78588 632120
rect 78088 632080 78588 632108
rect 78088 632068 78094 632080
rect 78582 632068 78588 632080
rect 78640 632068 78646 632120
rect 108942 632068 108948 632120
rect 109000 632108 109006 632120
rect 111794 632108 111800 632120
rect 109000 632080 111800 632108
rect 109000 632068 109006 632080
rect 111794 632068 111800 632080
rect 111852 632068 111858 632120
rect 115842 632068 115848 632120
rect 115900 632108 115906 632120
rect 121546 632108 121552 632120
rect 115900 632080 121552 632108
rect 115900 632068 115906 632080
rect 121546 632068 121552 632080
rect 121604 632068 121610 632120
rect 237926 632068 237932 632120
rect 237984 632108 237990 632120
rect 238662 632108 238668 632120
rect 237984 632080 238668 632108
rect 237984 632068 237990 632080
rect 238662 632068 238668 632080
rect 238720 632068 238726 632120
rect 255314 632068 255320 632120
rect 255372 632108 255378 632120
rect 256878 632108 256884 632120
rect 255372 632080 256884 632108
rect 255372 632068 255378 632080
rect 256878 632068 256884 632080
rect 256936 632068 256942 632120
rect 259362 632068 259368 632120
rect 259420 632108 259426 632120
rect 261754 632108 261760 632120
rect 259420 632080 261760 632108
rect 259420 632068 259426 632080
rect 261754 632068 261760 632080
rect 261812 632068 261818 632120
rect 482002 632068 482008 632120
rect 482060 632108 482066 632120
rect 482922 632108 482928 632120
rect 482060 632080 482928 632108
rect 482060 632068 482066 632080
rect 482922 632068 482928 632080
rect 482980 632068 482986 632120
rect 491846 632068 491852 632120
rect 491904 632108 491910 632120
rect 493318 632108 493324 632120
rect 491904 632080 493324 632108
rect 491904 632068 491910 632080
rect 493318 632068 493324 632080
rect 493376 632068 493382 632120
rect 500218 632068 500224 632120
rect 500276 632108 500282 632120
rect 501598 632108 501604 632120
rect 500276 632080 501604 632108
rect 500276 632068 500282 632080
rect 501598 632068 501604 632080
rect 501656 632068 501662 632120
rect 538858 630640 538864 630692
rect 538916 630680 538922 630692
rect 580166 630680 580172 630692
rect 538916 630652 580172 630680
rect 538916 630640 538922 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 72786 628260 72792 628312
rect 72844 628300 72850 628312
rect 232866 628300 232872 628312
rect 72844 628272 232872 628300
rect 72844 628260 72850 628272
rect 232866 628260 232872 628272
rect 232924 628260 232930 628312
rect 72694 628192 72700 628244
rect 72752 628232 72758 628244
rect 130378 628232 130384 628244
rect 72752 628204 130384 628232
rect 72752 628192 72758 628204
rect 130378 628192 130384 628204
rect 130436 628192 130442 628244
rect 232682 628192 232688 628244
rect 232740 628232 232746 628244
rect 289262 628232 289268 628244
rect 232740 628204 289268 628232
rect 232740 628192 232746 628204
rect 289262 628192 289268 628204
rect 289320 628192 289326 628244
rect 73062 628124 73068 628176
rect 73120 628164 73126 628176
rect 130562 628164 130568 628176
rect 73120 628136 130568 628164
rect 73120 628124 73126 628136
rect 130562 628124 130568 628136
rect 130620 628124 130626 628176
rect 233142 628124 233148 628176
rect 233200 628164 233206 628176
rect 290366 628164 290372 628176
rect 233200 628136 290372 628164
rect 233200 628124 233206 628136
rect 290366 628124 290372 628136
rect 290424 628124 290430 628176
rect 72602 628056 72608 628108
rect 72660 628096 72666 628108
rect 133138 628096 133144 628108
rect 72660 628068 133144 628096
rect 72660 628056 72666 628068
rect 133138 628056 133144 628068
rect 133196 628056 133202 628108
rect 235258 628056 235264 628108
rect 235316 628096 235322 628108
rect 290458 628096 290464 628108
rect 235316 628068 290464 628096
rect 235316 628056 235322 628068
rect 290458 628056 290464 628068
rect 290516 628056 290522 628108
rect 74442 627988 74448 628040
rect 74500 628028 74506 628040
rect 74500 628000 135208 628028
rect 74500 627988 74506 628000
rect 135180 627892 135208 628000
rect 232866 627988 232872 628040
rect 232924 628028 232930 628040
rect 313918 628028 313924 628040
rect 232924 628000 313924 628028
rect 232924 627988 232930 628000
rect 313918 627988 313924 628000
rect 313976 627988 313982 628040
rect 232774 627920 232780 627972
rect 232832 627960 232838 627972
rect 320818 627960 320824 627972
rect 232832 627932 320824 627960
rect 232832 627920 232838 627932
rect 320818 627920 320824 627932
rect 320876 627920 320882 627972
rect 233142 627892 233148 627904
rect 135180 627864 233148 627892
rect 233142 627852 233148 627864
rect 233200 627852 233206 627904
rect 72970 627648 72976 627700
rect 73028 627688 73034 627700
rect 128998 627688 129004 627700
rect 73028 627660 129004 627688
rect 73028 627648 73034 627660
rect 128998 627648 129004 627660
rect 129056 627648 129062 627700
rect 233050 627648 233056 627700
rect 233108 627688 233114 627700
rect 289078 627688 289084 627700
rect 233108 627660 289084 627688
rect 233108 627648 233114 627660
rect 289078 627648 289084 627660
rect 289136 627648 289142 627700
rect 72878 627580 72884 627632
rect 72936 627620 72942 627632
rect 130470 627620 130476 627632
rect 72936 627592 130476 627620
rect 72936 627580 72942 627592
rect 130470 627580 130476 627592
rect 130528 627580 130534 627632
rect 232958 627580 232964 627632
rect 233016 627620 233022 627632
rect 289170 627620 289176 627632
rect 233016 627592 289176 627620
rect 233016 627580 233022 627592
rect 289170 627580 289176 627592
rect 289228 627580 289234 627632
rect 290458 627172 290464 627224
rect 290516 627212 290522 627224
rect 454034 627212 454040 627224
rect 290516 627184 454040 627212
rect 290516 627172 290522 627184
rect 454034 627172 454040 627184
rect 454092 627172 454098 627224
rect 454034 626560 454040 626612
rect 454092 626600 454098 626612
rect 472618 626600 472624 626612
rect 454092 626572 472624 626600
rect 454092 626560 454098 626572
rect 472618 626560 472624 626572
rect 472676 626560 472682 626612
rect 133138 623704 133144 623756
rect 133196 623744 133202 623756
rect 232774 623744 232780 623756
rect 133196 623716 232780 623744
rect 133196 623704 133202 623716
rect 232774 623704 232780 623716
rect 232832 623704 232838 623756
rect 320818 623024 320824 623076
rect 320876 623064 320882 623076
rect 472158 623064 472164 623076
rect 320876 623036 472164 623064
rect 320876 623024 320882 623036
rect 472158 623024 472164 623036
rect 472216 623064 472222 623076
rect 472526 623064 472532 623076
rect 472216 623036 472532 623064
rect 472216 623024 472222 623036
rect 472526 623024 472532 623036
rect 472584 623024 472590 623076
rect 130562 619556 130568 619608
rect 130620 619596 130626 619608
rect 232314 619596 232320 619608
rect 130620 619568 232320 619596
rect 130620 619556 130626 619568
rect 232314 619556 232320 619568
rect 232372 619556 232378 619608
rect 289262 618876 289268 618928
rect 289320 618916 289326 618928
rect 451274 618916 451280 618928
rect 289320 618888 451280 618916
rect 289320 618876 289326 618888
rect 451274 618876 451280 618888
rect 451332 618916 451338 618928
rect 452194 618916 452200 618928
rect 451332 618888 452200 618916
rect 451332 618876 451338 618888
rect 452194 618876 452200 618888
rect 452252 618876 452258 618928
rect 452194 618264 452200 618316
rect 452252 618304 452258 618316
rect 472618 618304 472624 618316
rect 452252 618276 472624 618304
rect 452252 618264 452258 618276
rect 472618 618264 472624 618276
rect 472676 618264 472682 618316
rect 313918 614728 313924 614780
rect 313976 614768 313982 614780
rect 472250 614768 472256 614780
rect 313976 614740 472256 614768
rect 313976 614728 313982 614740
rect 472250 614728 472256 614740
rect 472308 614768 472314 614780
rect 472526 614768 472532 614780
rect 472308 614740 472532 614768
rect 472308 614728 472314 614740
rect 472526 614728 472532 614740
rect 472584 614728 472590 614780
rect 130470 611260 130476 611312
rect 130528 611300 130534 611312
rect 232958 611300 232964 611312
rect 130528 611272 232964 611300
rect 130528 611260 130534 611272
rect 232958 611260 232964 611272
rect 233016 611260 233022 611312
rect 289170 610580 289176 610632
rect 289228 610620 289234 610632
rect 449894 610620 449900 610632
rect 289228 610592 449900 610620
rect 289228 610580 289234 610592
rect 449894 610580 449900 610592
rect 449952 610580 449958 610632
rect 449894 609968 449900 610020
rect 449952 610008 449958 610020
rect 472618 610008 472624 610020
rect 449952 609980 472624 610008
rect 449952 609968 449958 609980
rect 472618 609968 472624 609980
rect 472676 609968 472682 610020
rect 128998 607112 129004 607164
rect 129056 607152 129062 607164
rect 232406 607152 232412 607164
rect 129056 607124 232412 607152
rect 129056 607112 129062 607124
rect 232406 607112 232412 607124
rect 232464 607112 232470 607164
rect 289078 606432 289084 606484
rect 289136 606472 289142 606484
rect 472434 606472 472440 606484
rect 289136 606444 472440 606472
rect 289136 606432 289142 606444
rect 472434 606432 472440 606444
rect 472492 606432 472498 606484
rect 130378 603032 130384 603084
rect 130436 603072 130442 603084
rect 233142 603072 233148 603084
rect 130436 603044 233148 603072
rect 130436 603032 130442 603044
rect 233142 603032 233148 603044
rect 233200 603032 233206 603084
rect 290458 602352 290464 602404
rect 290516 602392 290522 602404
rect 447134 602392 447140 602404
rect 290516 602364 447140 602392
rect 290516 602352 290522 602364
rect 447134 602352 447140 602364
rect 447192 602352 447198 602404
rect 447134 601672 447140 601724
rect 447192 601712 447198 601724
rect 472618 601712 472624 601724
rect 447192 601684 472624 601712
rect 447192 601672 447198 601684
rect 472618 601672 472624 601684
rect 472676 601672 472682 601724
rect 445018 589296 445024 589348
rect 445076 589336 445082 589348
rect 472618 589336 472624 589348
rect 445076 589308 472624 589336
rect 445076 589296 445082 589308
rect 472618 589296 472624 589308
rect 472676 589296 472682 589348
rect 459462 585148 459468 585200
rect 459520 585188 459526 585200
rect 472618 585188 472624 585200
rect 459520 585160 472624 585188
rect 459520 585148 459526 585160
rect 472618 585148 472624 585160
rect 472676 585148 472682 585200
rect 72786 582224 72792 582276
rect 72844 582264 72850 582276
rect 72970 582264 72976 582276
rect 72844 582236 72976 582264
rect 72844 582224 72850 582236
rect 72970 582224 72976 582236
rect 73028 582224 73034 582276
rect 444374 578144 444380 578196
rect 444432 578184 444438 578196
rect 445018 578184 445024 578196
rect 444432 578156 445024 578184
rect 444432 578144 444438 578156
rect 445018 578144 445024 578156
rect 445076 578144 445082 578196
rect 472526 578144 472532 578196
rect 472584 578184 472590 578196
rect 472986 578184 472992 578196
rect 472584 578156 472992 578184
rect 472584 578144 472590 578156
rect 472986 578144 472992 578156
rect 473044 578144 473050 578196
rect 472434 578076 472440 578128
rect 472492 578116 472498 578128
rect 473078 578116 473084 578128
rect 472492 578088 473084 578116
rect 472492 578076 472498 578088
rect 473078 578076 473084 578088
rect 473136 578076 473142 578128
rect 472526 577844 472532 577856
rect 451246 577816 472532 577844
rect 231762 577736 231768 577788
rect 231820 577776 231826 577788
rect 451246 577776 451274 577816
rect 472526 577804 472532 577816
rect 472584 577804 472590 577856
rect 231820 577748 451274 577776
rect 231820 577736 231826 577748
rect 72878 577668 72884 577720
rect 72936 577708 72942 577720
rect 232958 577708 232964 577720
rect 72936 577680 232964 577708
rect 72936 577668 72942 577680
rect 232958 577668 232964 577680
rect 233016 577708 233022 577720
rect 233016 577680 451274 577708
rect 233016 577668 233022 577680
rect 72970 577600 72976 577652
rect 73028 577640 73034 577652
rect 232774 577640 232780 577652
rect 73028 577612 232780 577640
rect 73028 577600 73034 577612
rect 232774 577600 232780 577612
rect 232832 577640 232838 577652
rect 444374 577640 444380 577652
rect 232832 577612 444380 577640
rect 232832 577600 232838 577612
rect 444374 577600 444380 577612
rect 444432 577600 444438 577652
rect 72786 577532 72792 577584
rect 72844 577572 72850 577584
rect 231762 577572 231768 577584
rect 72844 577544 231768 577572
rect 72844 577532 72850 577544
rect 231762 577532 231768 577544
rect 231820 577532 231826 577584
rect 451246 577572 451274 577680
rect 472434 577572 472440 577584
rect 451246 577544 472440 577572
rect 472434 577532 472440 577544
rect 472492 577532 472498 577584
rect 75822 577464 75828 577516
rect 75880 577504 75886 577516
rect 233142 577504 233148 577516
rect 75880 577476 233148 577504
rect 75880 577464 75886 577476
rect 233142 577464 233148 577476
rect 233200 577464 233206 577516
rect 235258 577464 235264 577516
rect 235316 577504 235322 577516
rect 472618 577504 472624 577516
rect 235316 577476 472624 577504
rect 235316 577464 235322 577476
rect 472618 577464 472624 577476
rect 472676 577464 472682 577516
rect 73062 577396 73068 577448
rect 73120 577436 73126 577448
rect 233050 577436 233056 577448
rect 73120 577408 233056 577436
rect 73120 577396 73126 577408
rect 233050 577396 233056 577408
rect 233108 577396 233114 577448
rect 17862 576852 17868 576904
rect 17920 576892 17926 576904
rect 71774 576892 71780 576904
rect 17920 576864 71780 576892
rect 17920 576852 17926 576864
rect 71774 576852 71780 576864
rect 71832 576852 71838 576904
rect 537478 576852 537484 576904
rect 537536 576892 537542 576904
rect 580166 576892 580172 576904
rect 537536 576864 580172 576892
rect 537536 576852 537542 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 233050 576172 233056 576224
rect 233108 576212 233114 576224
rect 339402 576212 339408 576224
rect 233108 576184 339408 576212
rect 233108 576172 233114 576184
rect 339402 576172 339408 576184
rect 339460 576172 339466 576224
rect 3510 576104 3516 576156
rect 3568 576144 3574 576156
rect 331858 576144 331864 576156
rect 3568 576116 331864 576144
rect 3568 576104 3574 576116
rect 331858 576104 331864 576116
rect 331916 576104 331922 576156
rect 475378 576104 475384 576156
rect 475436 576104 475442 576156
rect 480162 576104 480168 576156
rect 480220 576144 480226 576156
rect 528554 576144 528560 576156
rect 480220 576116 528560 576144
rect 480220 576104 480226 576116
rect 528554 576104 528560 576116
rect 528612 576104 528618 576156
rect 475396 575884 475424 576104
rect 475378 575832 475384 575884
rect 475436 575832 475442 575884
rect 339402 575424 339408 575476
rect 339460 575464 339466 575476
rect 473170 575464 473176 575476
rect 339460 575436 473176 575464
rect 339460 575424 339466 575436
rect 473170 575424 473176 575436
rect 473228 575424 473234 575476
rect 86126 573996 86132 574048
rect 86184 574036 86190 574048
rect 360286 574036 360292 574048
rect 86184 574008 360292 574036
rect 86184 573996 86190 574008
rect 360286 573996 360292 574008
rect 360344 573996 360350 574048
rect 426342 573996 426348 574048
rect 426400 574036 426406 574048
rect 519630 574036 519636 574048
rect 426400 574008 519636 574036
rect 426400 573996 426406 574008
rect 519630 573996 519636 574008
rect 519688 573996 519694 574048
rect 76374 573928 76380 573980
rect 76432 573968 76438 573980
rect 351914 573968 351920 573980
rect 76432 573940 351920 573968
rect 76432 573928 76438 573940
rect 351914 573928 351920 573940
rect 351972 573928 351978 573980
rect 367002 573928 367008 573980
rect 367060 573968 367066 573980
rect 488534 573968 488540 573980
rect 367060 573940 488540 573968
rect 367060 573928 367066 573940
rect 488534 573928 488540 573940
rect 488592 573928 488598 573980
rect 89438 573860 89444 573912
rect 89496 573900 89502 573912
rect 367094 573900 367100 573912
rect 89496 573872 367100 573900
rect 89496 573860 89502 573872
rect 367094 573860 367100 573872
rect 367152 573860 367158 573912
rect 369762 573860 369768 573912
rect 369820 573900 369826 573912
rect 490190 573900 490196 573912
rect 369820 573872 490196 573900
rect 369820 573860 369826 573872
rect 490190 573860 490196 573872
rect 490248 573860 490254 573912
rect 114002 573792 114008 573844
rect 114060 573832 114066 573844
rect 395338 573832 395344 573844
rect 114060 573804 395344 573832
rect 114060 573792 114066 573804
rect 395338 573792 395344 573804
rect 395396 573792 395402 573844
rect 407022 573792 407028 573844
rect 407080 573832 407086 573844
rect 509786 573832 509792 573844
rect 407080 573804 509792 573832
rect 407080 573792 407086 573804
rect 509786 573792 509792 573804
rect 509844 573792 509850 573844
rect 112346 573724 112352 573776
rect 112404 573764 112410 573776
rect 399478 573764 399484 573776
rect 112404 573736 399484 573764
rect 112404 573724 112410 573736
rect 399478 573724 399484 573736
rect 399536 573724 399542 573776
rect 404262 573724 404268 573776
rect 404320 573764 404326 573776
rect 508130 573764 508136 573776
rect 404320 573736 508136 573764
rect 404320 573724 404326 573736
rect 508130 573724 508136 573736
rect 508188 573724 508194 573776
rect 120534 573656 120540 573708
rect 120592 573696 120598 573708
rect 410518 573696 410524 573708
rect 120592 573668 410524 573696
rect 120592 573656 120598 573668
rect 410518 573656 410524 573668
rect 410576 573656 410582 573708
rect 416682 573656 416688 573708
rect 416740 573696 416746 573708
rect 514662 573696 514668 573708
rect 416740 573668 514668 573696
rect 416740 573656 416746 573668
rect 514662 573656 514668 573668
rect 514720 573656 514726 573708
rect 117222 573588 117228 573640
rect 117280 573628 117286 573640
rect 407758 573628 407764 573640
rect 117280 573600 407764 573628
rect 117280 573588 117286 573600
rect 407758 573588 407764 573600
rect 407816 573588 407822 573640
rect 411898 573588 411904 573640
rect 411956 573628 411962 573640
rect 511442 573628 511448 573640
rect 411956 573600 511448 573628
rect 411956 573588 411962 573600
rect 511442 573588 511448 573600
rect 511500 573588 511506 573640
rect 122190 573520 122196 573572
rect 122248 573560 122254 573572
rect 417418 573560 417424 573572
rect 122248 573532 417424 573560
rect 122248 573520 122254 573532
rect 417418 573520 417424 573532
rect 417476 573520 417482 573572
rect 419442 573520 419448 573572
rect 419500 573560 419506 573572
rect 516318 573560 516324 573572
rect 419500 573532 516324 573560
rect 419500 573520 419506 573532
rect 516318 573520 516324 573532
rect 516376 573520 516382 573572
rect 118510 573452 118516 573504
rect 118568 573492 118574 573504
rect 413278 573492 413284 573504
rect 118568 573464 413284 573492
rect 118568 573452 118574 573464
rect 413278 573452 413284 573464
rect 413336 573452 413342 573504
rect 414658 573452 414664 573504
rect 414716 573492 414722 573504
rect 513098 573492 513104 573504
rect 414716 573464 513104 573492
rect 414716 573452 414722 573464
rect 513098 573452 513104 573464
rect 513156 573452 513162 573504
rect 123754 573384 123760 573436
rect 123812 573424 123818 573436
rect 421558 573424 421564 573436
rect 123812 573396 421564 573424
rect 123812 573384 123818 573396
rect 421558 573384 421564 573396
rect 421616 573384 421622 573436
rect 423582 573384 423588 573436
rect 423640 573424 423646 573436
rect 517974 573424 517980 573436
rect 423640 573396 517980 573424
rect 423640 573384 423646 573396
rect 517974 573384 517980 573396
rect 518032 573384 518038 573436
rect 125410 573316 125416 573368
rect 125468 573356 125474 573368
rect 431218 573356 431224 573368
rect 125468 573328 431224 573356
rect 125468 573316 125474 573328
rect 431218 573316 431224 573328
rect 431276 573316 431282 573368
rect 433242 573316 433248 573368
rect 433300 573356 433306 573368
rect 522850 573356 522856 573368
rect 433300 573328 522856 573356
rect 433300 573316 433306 573328
rect 522850 573316 522856 573328
rect 522908 573316 522914 573368
rect 84102 573248 84108 573300
rect 84160 573288 84166 573300
rect 357434 573288 357440 573300
rect 84160 573260 357440 573288
rect 84160 573248 84166 573260
rect 357434 573248 357440 573260
rect 357492 573248 357498 573300
rect 429102 573248 429108 573300
rect 429160 573288 429166 573300
rect 521286 573288 521292 573300
rect 429160 573260 521292 573288
rect 429160 573248 429166 573260
rect 521286 573248 521292 573260
rect 521344 573248 521350 573300
rect 87782 573180 87788 573232
rect 87840 573220 87846 573232
rect 98641 573223 98699 573229
rect 98641 573220 98653 573223
rect 87840 573192 98653 573220
rect 87840 573180 87846 573192
rect 98641 573189 98653 573192
rect 98687 573189 98699 573223
rect 98641 573183 98699 573189
rect 104158 573180 104164 573232
rect 104216 573220 104222 573232
rect 106918 573220 106924 573232
rect 104216 573192 106924 573220
rect 104216 573180 104222 573192
rect 106918 573180 106924 573192
rect 106976 573180 106982 573232
rect 115566 573180 115572 573232
rect 115624 573220 115630 573232
rect 363598 573220 363604 573232
rect 115624 573192 363604 573220
rect 115624 573180 115630 573192
rect 363598 573180 363604 573192
rect 363656 573180 363662 573232
rect 436002 573180 436008 573232
rect 436060 573220 436066 573232
rect 524506 573220 524512 573232
rect 436060 573192 524512 573220
rect 436060 573180 436066 573192
rect 524506 573180 524512 573192
rect 524564 573180 524570 573232
rect 82722 573112 82728 573164
rect 82780 573152 82786 573164
rect 327718 573152 327724 573164
rect 82780 573124 327724 573152
rect 82780 573112 82786 573124
rect 327718 573112 327724 573124
rect 327776 573112 327782 573164
rect 438762 573112 438768 573164
rect 438820 573152 438826 573164
rect 526162 573152 526168 573164
rect 438820 573124 526168 573152
rect 438820 573112 438826 573124
rect 526162 573112 526168 573124
rect 526220 573112 526226 573164
rect 98641 573087 98699 573093
rect 98641 573053 98653 573087
rect 98687 573084 98699 573087
rect 331950 573084 331956 573096
rect 98687 573056 331956 573084
rect 98687 573053 98699 573056
rect 98641 573047 98699 573053
rect 331950 573044 331956 573056
rect 332008 573044 332014 573096
rect 441522 573044 441528 573096
rect 441580 573084 441586 573096
rect 527818 573084 527824 573096
rect 441580 573056 527824 573084
rect 441580 573044 441586 573056
rect 527818 573044 527824 573056
rect 527876 573044 527882 573096
rect 91002 572976 91008 573028
rect 91060 573016 91066 573028
rect 334710 573016 334716 573028
rect 91060 572988 334716 573016
rect 91060 572976 91066 572988
rect 334710 572976 334716 572988
rect 334768 572976 334774 573028
rect 409138 572976 409144 573028
rect 409196 573016 409202 573028
rect 478690 573016 478696 573028
rect 409196 572988 478696 573016
rect 409196 572976 409202 572988
rect 478690 572976 478696 572988
rect 478748 572976 478754 573028
rect 482278 572976 482284 573028
rect 482336 573016 482342 573028
rect 491754 573016 491760 573028
rect 482336 572988 491760 573016
rect 482336 572976 482342 572988
rect 491754 572976 491760 572988
rect 491812 572976 491818 573028
rect 81250 572908 81256 572960
rect 81308 572948 81314 572960
rect 322198 572948 322204 572960
rect 81308 572920 322204 572948
rect 81308 572908 81314 572920
rect 322198 572908 322204 572920
rect 322256 572908 322262 572960
rect 420178 572908 420184 572960
rect 420236 572948 420242 572960
rect 480346 572948 480352 572960
rect 420236 572920 480352 572948
rect 420236 572908 420242 572920
rect 480346 572908 480352 572920
rect 480404 572908 480410 572960
rect 480809 572951 480867 572957
rect 480809 572917 480821 572951
rect 480855 572948 480867 572951
rect 485222 572948 485228 572960
rect 480855 572920 485228 572948
rect 480855 572917 480867 572920
rect 480809 572911 480867 572917
rect 485222 572908 485228 572920
rect 485280 572908 485286 572960
rect 102502 572840 102508 572892
rect 102560 572880 102566 572892
rect 105538 572880 105544 572892
rect 102560 572852 105544 572880
rect 102560 572840 102566 572852
rect 105538 572840 105544 572852
rect 105596 572840 105602 572892
rect 126882 572840 126888 572892
rect 126940 572880 126946 572892
rect 323578 572880 323584 572892
rect 126940 572852 323584 572880
rect 126940 572840 126946 572852
rect 323578 572840 323584 572852
rect 323636 572840 323642 572892
rect 443638 572840 443644 572892
rect 443696 572880 443702 572892
rect 482002 572880 482008 572892
rect 443696 572852 482008 572880
rect 443696 572840 443702 572852
rect 482002 572840 482008 572852
rect 482060 572840 482066 572892
rect 100662 572772 100668 572824
rect 100720 572812 100726 572824
rect 104158 572812 104164 572824
rect 100720 572784 104164 572812
rect 100720 572772 100726 572784
rect 104158 572772 104164 572784
rect 104216 572772 104222 572824
rect 128722 572772 128728 572824
rect 128780 572812 128786 572824
rect 324958 572812 324964 572824
rect 128780 572784 324964 572812
rect 128780 572772 128786 572784
rect 324958 572772 324964 572784
rect 325016 572772 325022 572824
rect 476758 572772 476764 572824
rect 476816 572812 476822 572824
rect 483566 572812 483572 572824
rect 476816 572784 483572 572812
rect 476816 572772 476822 572784
rect 483566 572772 483572 572784
rect 483624 572772 483630 572824
rect 77938 572704 77944 572756
rect 77996 572744 78002 572756
rect 78582 572744 78588 572756
rect 77996 572716 78588 572744
rect 77996 572704 78002 572716
rect 78582 572704 78588 572716
rect 78640 572704 78646 572756
rect 94314 572704 94320 572756
rect 94372 572744 94378 572756
rect 95142 572744 95148 572756
rect 94372 572716 95148 572744
rect 94372 572704 94378 572716
rect 95142 572704 95148 572716
rect 95200 572704 95206 572756
rect 95970 572704 95976 572756
rect 96028 572744 96034 572756
rect 97258 572744 97264 572756
rect 96028 572716 97264 572744
rect 96028 572704 96034 572716
rect 97258 572704 97264 572716
rect 97316 572704 97322 572756
rect 97626 572704 97632 572756
rect 97684 572744 97690 572756
rect 98638 572744 98644 572756
rect 97684 572716 98644 572744
rect 97684 572704 97690 572716
rect 98638 572704 98644 572716
rect 98696 572704 98702 572756
rect 99282 572704 99288 572756
rect 99340 572744 99346 572756
rect 101398 572744 101404 572756
rect 99340 572716 101404 572744
rect 99340 572704 99346 572716
rect 101398 572704 101404 572716
rect 101456 572704 101462 572756
rect 105814 572704 105820 572756
rect 105872 572744 105878 572756
rect 108298 572744 108304 572756
rect 105872 572716 108304 572744
rect 105872 572704 105878 572716
rect 108298 572704 108304 572716
rect 108356 572704 108362 572756
rect 108942 572704 108948 572756
rect 109000 572744 109006 572756
rect 111058 572744 111064 572756
rect 109000 572716 111064 572744
rect 109000 572704 109006 572716
rect 111058 572704 111064 572716
rect 111116 572704 111122 572756
rect 237834 572704 237840 572756
rect 237892 572744 237898 572756
rect 238662 572744 238668 572756
rect 237892 572716 238668 572744
rect 237892 572704 237898 572716
rect 238662 572704 238668 572716
rect 238720 572704 238726 572756
rect 246022 572704 246028 572756
rect 246080 572744 246086 572756
rect 246942 572744 246948 572756
rect 246080 572716 246948 572744
rect 246080 572704 246086 572716
rect 246942 572704 246948 572716
rect 247000 572704 247006 572756
rect 255866 572704 255872 572756
rect 255924 572744 255930 572756
rect 256602 572744 256608 572756
rect 255924 572716 256608 572744
rect 255924 572704 255930 572716
rect 256602 572704 256608 572716
rect 256660 572704 256666 572756
rect 264054 572704 264060 572756
rect 264112 572744 264118 572756
rect 264882 572744 264888 572756
rect 264112 572716 264888 572744
rect 264112 572704 264118 572716
rect 264882 572704 264888 572716
rect 264940 572704 264946 572756
rect 272242 572704 272248 572756
rect 272300 572744 272306 572756
rect 273162 572744 273168 572756
rect 272300 572716 273168 572744
rect 272300 572704 272306 572716
rect 273162 572704 273168 572716
rect 273220 572704 273226 572756
rect 273898 572704 273904 572756
rect 273956 572744 273962 572756
rect 274542 572744 274548 572756
rect 273956 572716 274548 572744
rect 273956 572704 273962 572716
rect 274542 572704 274548 572716
rect 274600 572704 274606 572756
rect 275462 572704 275468 572756
rect 275520 572744 275526 572756
rect 275922 572744 275928 572756
rect 275520 572716 275928 572744
rect 275520 572704 275526 572716
rect 275922 572704 275928 572716
rect 275980 572704 275986 572756
rect 280430 572704 280436 572756
rect 280488 572744 280494 572756
rect 281442 572744 281448 572756
rect 280488 572716 281448 572744
rect 280488 572704 280494 572716
rect 281442 572704 281448 572716
rect 281500 572704 281506 572756
rect 282086 572704 282092 572756
rect 282144 572744 282150 572756
rect 282822 572744 282828 572756
rect 282144 572716 282828 572744
rect 282144 572704 282150 572716
rect 282822 572704 282828 572716
rect 282880 572704 282886 572756
rect 283650 572704 283656 572756
rect 283708 572744 283714 572756
rect 284202 572744 284208 572756
rect 283708 572716 284208 572744
rect 283708 572704 283714 572716
rect 284202 572704 284208 572716
rect 284260 572704 284266 572756
rect 478138 572704 478144 572756
rect 478196 572744 478202 572756
rect 480809 572747 480867 572753
rect 480809 572744 480821 572747
rect 478196 572716 480821 572744
rect 478196 572704 478202 572716
rect 480809 572713 480821 572716
rect 480855 572713 480867 572747
rect 480809 572707 480867 572713
rect 480898 572704 480904 572756
rect 480956 572744 480962 572756
rect 486878 572744 486884 572756
rect 480956 572716 486884 572744
rect 480956 572704 480962 572716
rect 486878 572704 486884 572716
rect 486936 572704 486942 572756
rect 497458 572704 497464 572756
rect 497516 572744 497522 572756
rect 498378 572744 498384 572756
rect 497516 572716 498384 572744
rect 497516 572704 497522 572716
rect 498378 572704 498384 572716
rect 498436 572704 498442 572756
rect 247678 572636 247684 572688
rect 247736 572676 247742 572688
rect 349798 572676 349804 572688
rect 247736 572648 349804 572676
rect 247736 572636 247742 572648
rect 349798 572636 349804 572648
rect 349856 572636 349862 572688
rect 236270 572568 236276 572620
rect 236328 572608 236334 572620
rect 341518 572608 341524 572620
rect 236328 572580 341524 572608
rect 236328 572568 236334 572580
rect 341518 572568 341524 572580
rect 341576 572568 341582 572620
rect 239490 572500 239496 572552
rect 239548 572540 239554 572552
rect 345014 572540 345020 572552
rect 239548 572512 345020 572540
rect 239548 572500 239554 572512
rect 345014 572500 345020 572512
rect 345072 572500 345078 572552
rect 244182 572432 244188 572484
rect 244240 572472 244246 572484
rect 356054 572472 356060 572484
rect 244240 572444 356060 572472
rect 244240 572432 244246 572444
rect 356054 572432 356060 572444
rect 356112 572432 356118 572484
rect 257522 572364 257528 572416
rect 257580 572404 257586 572416
rect 370498 572404 370504 572416
rect 257580 572376 370504 572404
rect 257580 572364 257586 572376
rect 370498 572364 370504 572376
rect 370556 572364 370562 572416
rect 382182 572364 382188 572416
rect 382240 572404 382246 572416
rect 496722 572404 496728 572416
rect 382240 572376 496728 572404
rect 382240 572364 382246 572376
rect 496722 572364 496728 572376
rect 496780 572364 496786 572416
rect 254210 572296 254216 572348
rect 254268 572336 254274 572348
rect 374638 572336 374644 572348
rect 254268 572308 374644 572336
rect 254268 572296 254274 572308
rect 374638 572296 374644 572308
rect 374696 572296 374702 572348
rect 379422 572296 379428 572348
rect 379480 572336 379486 572348
rect 495066 572336 495072 572348
rect 379480 572308 495072 572336
rect 379480 572296 379486 572308
rect 495066 572296 495072 572308
rect 495124 572296 495130 572348
rect 262122 572228 262128 572280
rect 262180 572268 262186 572280
rect 388438 572268 388444 572280
rect 262180 572240 388444 572268
rect 262180 572228 262186 572240
rect 388438 572228 388444 572240
rect 388496 572228 388502 572280
rect 265710 572160 265716 572212
rect 265768 572200 265774 572212
rect 396718 572200 396724 572212
rect 265768 572172 396724 572200
rect 265768 572160 265774 572172
rect 396718 572160 396724 572172
rect 396776 572160 396782 572212
rect 340782 572092 340788 572144
rect 340840 572132 340846 572144
rect 477034 572132 477040 572144
rect 340840 572104 477040 572132
rect 340840 572092 340846 572104
rect 477034 572092 477040 572104
rect 477092 572092 477098 572144
rect 110322 572024 110328 572076
rect 110380 572064 110386 572076
rect 382918 572064 382924 572076
rect 110380 572036 382924 572064
rect 110380 572024 110386 572036
rect 382918 572024 382924 572036
rect 382976 572024 382982 572076
rect 107378 571956 107384 572008
rect 107436 571996 107442 572008
rect 393958 571996 393964 572008
rect 107436 571968 393964 571996
rect 107436 571956 107442 571968
rect 393958 571956 393964 571968
rect 394016 571956 394022 572008
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 334618 565876 334624 565888
rect 3292 565848 334624 565876
rect 3292 565836 3298 565848
rect 334618 565836 334624 565848
rect 334676 565836 334682 565888
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 322290 553432 322296 553444
rect 3384 553404 322296 553432
rect 3384 553392 3390 553404
rect 322290 553392 322296 553404
rect 322348 553392 322354 553444
rect 482370 536800 482376 536852
rect 482428 536840 482434 536852
rect 579890 536840 579896 536852
rect 482428 536812 579896 536840
rect 482428 536800 482434 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 482462 524424 482468 524476
rect 482520 524464 482526 524476
rect 580166 524464 580172 524476
rect 482520 524436 580172 524464
rect 482520 524424 482526 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 500964 3516 501016
rect 3568 501004 3574 501016
rect 320910 501004 320916 501016
rect 3568 500976 320916 501004
rect 3568 500964 3574 500976
rect 320910 500964 320916 500976
rect 320968 500964 320974 501016
rect 482554 484372 482560 484424
rect 482612 484412 482618 484424
rect 580166 484412 580172 484424
rect 482612 484384 580172 484412
rect 482612 484372 482618 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 482646 470568 482652 470620
rect 482704 470608 482710 470620
rect 580166 470608 580172 470620
rect 482704 470580 580172 470608
rect 482704 470568 482710 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 330570 462380 330576 462392
rect 3568 462352 330576 462380
rect 3568 462340 3574 462352
rect 330570 462340 330576 462352
rect 330628 462340 330634 462392
rect 246942 456152 246948 456204
rect 247000 456192 247006 456204
rect 353938 456192 353944 456204
rect 247000 456164 353944 456192
rect 247000 456152 247006 456164
rect 353938 456152 353944 456164
rect 353996 456152 354002 456204
rect 260742 456084 260748 456136
rect 260800 456124 260806 456136
rect 387794 456124 387800 456136
rect 260800 456096 387800 456124
rect 260800 456084 260806 456096
rect 387794 456084 387800 456096
rect 387852 456084 387858 456136
rect 267642 456016 267648 456068
rect 267700 456056 267706 456068
rect 400214 456056 400220 456068
rect 267700 456028 400220 456056
rect 267700 456016 267706 456028
rect 400214 456016 400220 456028
rect 400272 456016 400278 456068
rect 238662 453364 238668 453416
rect 238720 453404 238726 453416
rect 340874 453404 340880 453416
rect 238720 453376 340880 453404
rect 238720 453364 238726 453376
rect 340874 453364 340880 453376
rect 340932 453364 340938 453416
rect 79962 453296 79968 453348
rect 80020 453336 80026 453348
rect 342898 453336 342904 453348
rect 80020 453308 342904 453336
rect 80020 453296 80026 453308
rect 342898 453296 342904 453308
rect 342956 453296 342962 453348
rect 3510 448536 3516 448588
rect 3568 448576 3574 448588
rect 325326 448576 325332 448588
rect 3568 448548 325332 448576
rect 3568 448536 3574 448548
rect 325326 448536 325332 448548
rect 325384 448536 325390 448588
rect 482738 430584 482744 430636
rect 482796 430624 482802 430636
rect 579890 430624 579896 430636
rect 482796 430596 579896 430624
rect 482796 430584 482802 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 482830 418140 482836 418192
rect 482888 418180 482894 418192
rect 580166 418180 580172 418192
rect 482888 418152 580172 418180
rect 482888 418140 482894 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 104158 412156 104164 412208
rect 104216 412196 104222 412208
rect 389450 412196 389456 412208
rect 104216 412168 389456 412196
rect 104216 412156 104222 412168
rect 389450 412156 389456 412168
rect 389508 412156 389514 412208
rect 105538 412088 105544 412140
rect 105596 412128 105602 412140
rect 392670 412128 392676 412140
rect 105596 412100 392676 412128
rect 105596 412088 105602 412100
rect 392670 412088 392676 412100
rect 392728 412088 392734 412140
rect 106918 412020 106924 412072
rect 106976 412060 106982 412072
rect 396074 412060 396080 412072
rect 106976 412032 396080 412060
rect 106976 412020 106982 412032
rect 396074 412020 396080 412032
rect 396132 412020 396138 412072
rect 108298 411952 108304 412004
rect 108356 411992 108362 412004
rect 398926 411992 398932 412004
rect 108356 411964 398932 411992
rect 108356 411952 108362 411964
rect 398926 411952 398932 411964
rect 398984 411952 398990 412004
rect 111058 411884 111064 411936
rect 111116 411924 111122 411936
rect 405734 411924 405740 411936
rect 111116 411896 405740 411924
rect 111116 411884 111122 411896
rect 405734 411884 405740 411896
rect 405792 411884 405798 411936
rect 251082 411204 251088 411256
rect 251140 411244 251146 411256
rect 369946 411244 369952 411256
rect 251140 411216 369952 411244
rect 251140 411204 251146 411216
rect 369946 411204 369952 411216
rect 370004 411204 370010 411256
rect 252462 411136 252468 411188
rect 252520 411176 252526 411188
rect 371878 411176 371884 411188
rect 252520 411148 371884 411176
rect 252520 411136 252526 411148
rect 371878 411136 371884 411148
rect 371936 411136 371942 411188
rect 256602 411068 256608 411120
rect 256660 411108 256666 411120
rect 378962 411108 378968 411120
rect 256660 411080 378968 411108
rect 256660 411068 256666 411080
rect 378962 411068 378968 411080
rect 379020 411068 379026 411120
rect 259362 411000 259368 411052
rect 259420 411040 259426 411052
rect 385310 411040 385316 411052
rect 259420 411012 385316 411040
rect 259420 411000 259426 411012
rect 385310 411000 385316 411012
rect 385368 411000 385374 411052
rect 264882 410932 264888 410984
rect 264940 410972 264946 410984
rect 394786 410972 394792 410984
rect 264940 410944 394792 410972
rect 264940 410932 264946 410944
rect 394786 410932 394792 410944
rect 394844 410932 394850 410984
rect 269022 410864 269028 410916
rect 269080 410904 269086 410916
rect 403618 410904 403624 410916
rect 269080 410876 403624 410904
rect 269080 410864 269086 410876
rect 403618 410864 403624 410876
rect 403676 410864 403682 410916
rect 273162 410796 273168 410848
rect 273220 410836 273226 410848
rect 410426 410836 410432 410848
rect 273220 410808 410432 410836
rect 273220 410796 273226 410808
rect 410426 410796 410432 410808
rect 410484 410796 410490 410848
rect 270402 410728 270408 410780
rect 270460 410768 270466 410780
rect 407390 410768 407396 410780
rect 270460 410740 407396 410768
rect 270460 410728 270466 410740
rect 407390 410728 407396 410740
rect 407448 410728 407454 410780
rect 274542 410660 274548 410712
rect 274600 410700 274606 410712
rect 414106 410700 414112 410712
rect 274600 410672 414112 410700
rect 274600 410660 274606 410672
rect 414106 410660 414112 410672
rect 414164 410660 414170 410712
rect 98638 410592 98644 410644
rect 98696 410632 98702 410644
rect 383654 410632 383660 410644
rect 98696 410604 383660 410632
rect 98696 410592 98702 410604
rect 383654 410592 383660 410604
rect 383712 410592 383718 410644
rect 101398 410524 101404 410576
rect 101456 410564 101462 410576
rect 386414 410564 386420 410576
rect 101456 410536 386420 410564
rect 101456 410524 101462 410536
rect 386414 410524 386420 410536
rect 386472 410524 386478 410576
rect 249702 410456 249708 410508
rect 249760 410496 249766 410508
rect 364978 410496 364984 410508
rect 249760 410468 364984 410496
rect 249760 410456 249766 410468
rect 364978 410456 364984 410468
rect 365036 410456 365042 410508
rect 228818 410184 228824 410236
rect 228876 410224 228882 410236
rect 327902 410224 327908 410236
rect 228876 410196 327908 410224
rect 228876 410184 228882 410196
rect 327902 410184 327908 410196
rect 327960 410184 327966 410236
rect 226242 410116 226248 410168
rect 226300 410156 226306 410168
rect 326338 410156 326344 410168
rect 226300 410128 326344 410156
rect 226300 410116 226306 410128
rect 326338 410116 326344 410128
rect 326396 410116 326402 410168
rect 222102 410048 222108 410100
rect 222160 410088 222166 410100
rect 325142 410088 325148 410100
rect 222160 410060 325148 410088
rect 222160 410048 222166 410060
rect 325142 410048 325148 410060
rect 325200 410048 325206 410100
rect 223482 409980 223488 410032
rect 223540 410020 223546 410032
rect 329190 410020 329196 410032
rect 223540 409992 329196 410020
rect 223540 409980 223546 409992
rect 329190 409980 329196 409992
rect 329248 409980 329254 410032
rect 218974 409912 218980 409964
rect 219032 409952 219038 409964
rect 332042 409952 332048 409964
rect 219032 409924 332048 409952
rect 219032 409912 219038 409924
rect 332042 409912 332048 409924
rect 332100 409912 332106 409964
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 329558 409884 329564 409896
rect 3200 409856 329564 409884
rect 3200 409844 3206 409856
rect 329558 409844 329564 409856
rect 329616 409844 329622 409896
rect 211062 409776 211068 409828
rect 211120 409816 211126 409828
rect 333238 409816 333244 409828
rect 211120 409788 333244 409816
rect 211120 409776 211126 409788
rect 333238 409776 333244 409788
rect 333296 409776 333302 409828
rect 3694 409708 3700 409760
rect 3752 409748 3758 409760
rect 328270 409748 328276 409760
rect 3752 409720 328276 409748
rect 3752 409708 3758 409720
rect 328270 409708 328276 409720
rect 328328 409708 328334 409760
rect 264882 409640 264888 409692
rect 264940 409680 264946 409692
rect 319530 409680 319536 409692
rect 264940 409652 319536 409680
rect 264940 409640 264946 409652
rect 319530 409640 319536 409652
rect 319588 409640 319594 409692
rect 278682 409572 278688 409624
rect 278740 409612 278746 409624
rect 337562 409612 337568 409624
rect 278740 409584 337568 409612
rect 278740 409572 278746 409584
rect 337562 409572 337568 409584
rect 337620 409572 337626 409624
rect 274542 409504 274548 409556
rect 274600 409544 274606 409556
rect 336550 409544 336556 409556
rect 274600 409516 336556 409544
rect 274600 409504 274606 409516
rect 336550 409504 336556 409516
rect 336608 409504 336614 409556
rect 271782 409436 271788 409488
rect 271840 409476 271846 409488
rect 335262 409476 335268 409488
rect 271840 409448 335268 409476
rect 271840 409436 271846 409448
rect 335262 409436 335268 409448
rect 335320 409436 335326 409488
rect 232866 409368 232872 409420
rect 232924 409408 232930 409420
rect 459002 409408 459008 409420
rect 232924 409380 459008 409408
rect 232924 409368 232930 409380
rect 459002 409368 459008 409380
rect 459060 409368 459066 409420
rect 78582 409300 78588 409352
rect 78640 409340 78646 409352
rect 342254 409340 342260 409352
rect 78640 409312 342260 409340
rect 78640 409300 78646 409312
rect 342254 409300 342260 409312
rect 342312 409300 342318 409352
rect 95142 409232 95148 409284
rect 95200 409272 95206 409284
rect 376846 409272 376852 409284
rect 95200 409244 376852 409272
rect 95200 409232 95206 409244
rect 376846 409232 376852 409244
rect 376904 409232 376910 409284
rect 92382 409164 92388 409216
rect 92440 409204 92446 409216
rect 373994 409204 374000 409216
rect 92440 409176 374000 409204
rect 92440 409164 92446 409176
rect 373994 409164 374000 409176
rect 374052 409164 374058 409216
rect 97258 409096 97264 409148
rect 97316 409136 97322 409148
rect 379974 409136 379980 409148
rect 97316 409108 379980 409136
rect 97316 409096 97322 409108
rect 379974 409096 379980 409108
rect 380032 409096 380038 409148
rect 259362 409028 259368 409080
rect 259420 409068 259426 409080
rect 326522 409068 326528 409080
rect 259420 409040 326528 409068
rect 259420 409028 259426 409040
rect 326522 409028 326528 409040
rect 326580 409028 326586 409080
rect 256602 408960 256608 409012
rect 256660 409000 256666 409012
rect 324038 409000 324044 409012
rect 256660 408972 324044 409000
rect 256660 408960 256666 408972
rect 324038 408960 324044 408972
rect 324096 408960 324102 409012
rect 266262 408892 266268 408944
rect 266320 408932 266326 408944
rect 337470 408932 337476 408944
rect 266320 408904 337476 408932
rect 266320 408892 266326 408904
rect 337470 408892 337476 408904
rect 337528 408892 337534 408944
rect 253842 408824 253848 408876
rect 253900 408864 253906 408876
rect 330754 408864 330760 408876
rect 253900 408836 330760 408864
rect 253900 408824 253906 408836
rect 330754 408824 330760 408836
rect 330812 408824 330818 408876
rect 251082 408756 251088 408808
rect 251140 408796 251146 408808
rect 329282 408796 329288 408808
rect 251140 408768 329288 408796
rect 251140 408756 251146 408768
rect 329282 408756 329288 408768
rect 329340 408756 329346 408808
rect 213822 408688 213828 408740
rect 213880 408728 213886 408740
rect 321002 408728 321008 408740
rect 213880 408700 321008 408728
rect 213880 408688 213886 408700
rect 321002 408688 321008 408700
rect 321060 408688 321066 408740
rect 216582 408620 216588 408672
rect 216640 408660 216646 408672
rect 337378 408660 337384 408672
rect 216640 408632 337384 408660
rect 216640 408620 216646 408632
rect 337378 408620 337384 408632
rect 337436 408620 337442 408672
rect 286502 408552 286508 408604
rect 286560 408592 286566 408604
rect 319438 408592 319444 408604
rect 286560 408564 319444 408592
rect 286560 408552 286566 408564
rect 319438 408552 319444 408564
rect 319496 408552 319502 408604
rect 276842 408484 276848 408536
rect 276900 408524 276906 408536
rect 322566 408524 322572 408536
rect 276900 408496 322572 408524
rect 276900 408484 276906 408496
rect 322566 408484 322572 408496
rect 322624 408484 322630 408536
rect 114462 408416 114468 408468
rect 114520 408456 114526 408468
rect 332410 408456 332416 408468
rect 114520 408428 332416 408456
rect 114520 408416 114526 408428
rect 332410 408416 332416 408428
rect 332468 408416 332474 408468
rect 124122 408348 124128 408400
rect 124180 408388 124186 408400
rect 318242 408388 318248 408400
rect 124180 408360 318248 408388
rect 124180 408348 124186 408360
rect 318242 408348 318248 408360
rect 318300 408348 318306 408400
rect 284202 408280 284208 408332
rect 284260 408320 284266 408332
rect 327994 408320 328000 408332
rect 284260 408292 328000 408320
rect 284260 408280 284266 408292
rect 327994 408280 328000 408292
rect 328052 408280 328058 408332
rect 269022 408212 269028 408264
rect 269080 408252 269086 408264
rect 318426 408252 318432 408264
rect 269080 408224 318432 408252
rect 269080 408212 269086 408224
rect 318426 408212 318432 408224
rect 318484 408212 318490 408264
rect 262122 408144 262128 408196
rect 262180 408184 262186 408196
rect 319622 408184 319628 408196
rect 262180 408156 319628 408184
rect 262180 408144 262186 408156
rect 319622 408144 319628 408156
rect 319680 408144 319686 408196
rect 249702 408076 249708 408128
rect 249760 408116 249766 408128
rect 325418 408116 325424 408128
rect 249760 408088 325424 408116
rect 249760 408076 249766 408088
rect 325418 408076 325424 408088
rect 325476 408076 325482 408128
rect 246942 408008 246948 408060
rect 247000 408048 247006 408060
rect 336274 408048 336280 408060
rect 247000 408020 336280 408048
rect 247000 408008 247006 408020
rect 336274 408008 336280 408020
rect 336332 408008 336338 408060
rect 140682 407940 140688 407992
rect 140740 407980 140746 407992
rect 157518 407980 157524 407992
rect 140740 407952 157524 407980
rect 140740 407940 140746 407952
rect 157518 407940 157524 407952
rect 157576 407940 157582 407992
rect 234522 407940 234528 407992
rect 234580 407980 234586 407992
rect 323854 407980 323860 407992
rect 234580 407952 323860 407980
rect 234580 407940 234586 407952
rect 323854 407940 323860 407952
rect 323912 407940 323918 407992
rect 139302 407872 139308 407924
rect 139360 407912 139366 407924
rect 157426 407912 157432 407924
rect 139360 407884 157432 407912
rect 139360 407872 139366 407884
rect 157426 407872 157432 407884
rect 157484 407872 157490 407924
rect 241422 407872 241428 407924
rect 241480 407912 241486 407924
rect 332226 407912 332232 407924
rect 241480 407884 332232 407912
rect 241480 407872 241486 407884
rect 332226 407872 332232 407884
rect 332284 407872 332290 407924
rect 71682 407804 71688 407856
rect 71740 407844 71746 407856
rect 156782 407844 156788 407856
rect 71740 407816 156788 407844
rect 71740 407804 71746 407816
rect 156782 407804 156788 407816
rect 156840 407804 156846 407856
rect 237282 407804 237288 407856
rect 237340 407844 237346 407856
rect 334894 407844 334900 407856
rect 237340 407816 334900 407844
rect 237340 407804 237346 407816
rect 334894 407804 334900 407816
rect 334952 407804 334958 407856
rect 66162 407736 66168 407788
rect 66220 407776 66226 407788
rect 156690 407776 156696 407788
rect 66220 407748 156696 407776
rect 66220 407736 66226 407748
rect 156690 407736 156696 407748
rect 156748 407736 156754 407788
rect 231762 407736 231768 407788
rect 231820 407776 231826 407788
rect 330846 407776 330852 407788
rect 231820 407748 330852 407776
rect 231820 407736 231826 407748
rect 330846 407736 330852 407748
rect 330904 407736 330910 407788
rect 64506 407668 64512 407720
rect 64564 407708 64570 407720
rect 156598 407708 156604 407720
rect 64564 407680 156604 407708
rect 64564 407668 64570 407680
rect 156598 407668 156604 407680
rect 156656 407668 156662 407720
rect 209498 407668 209504 407720
rect 209556 407708 209562 407720
rect 327810 407708 327816 407720
rect 209556 407680 327816 407708
rect 209556 407668 209562 407680
rect 327810 407668 327816 407680
rect 327868 407668 327874 407720
rect 121362 407600 121368 407652
rect 121420 407640 121426 407652
rect 322658 407640 322664 407652
rect 121420 407612 322664 407640
rect 121420 407600 121426 407612
rect 322658 407600 322664 407612
rect 322716 407600 322722 407652
rect 117222 407532 117228 407584
rect 117280 407572 117286 407584
rect 318518 407572 318524 407584
rect 117280 407544 318524 407572
rect 117280 407532 117286 407544
rect 318518 407532 318524 407544
rect 318576 407532 318582 407584
rect 126882 407464 126888 407516
rect 126940 407504 126946 407516
rect 329466 407504 329472 407516
rect 126940 407476 329472 407504
rect 126940 407464 126946 407476
rect 329466 407464 329472 407476
rect 329524 407464 329530 407516
rect 118602 407396 118608 407448
rect 118660 407436 118666 407448
rect 321370 407436 321376 407448
rect 118660 407408 321376 407436
rect 118660 407396 118666 407408
rect 321370 407396 321376 407408
rect 321428 407396 321434 407448
rect 111702 407328 111708 407380
rect 111760 407368 111766 407380
rect 328178 407368 328184 407380
rect 111760 407340 328184 407368
rect 111760 407328 111766 407340
rect 328178 407328 328184 407340
rect 328236 407328 328242 407380
rect 108942 407260 108948 407312
rect 109000 407300 109006 407312
rect 325510 407300 325516 407312
rect 109000 407272 325516 407300
rect 109000 407260 109006 407272
rect 325510 407260 325516 407272
rect 325568 407260 325574 407312
rect 300762 407192 300768 407244
rect 300820 407232 300826 407244
rect 317598 407232 317604 407244
rect 300820 407204 317604 407232
rect 300820 407192 300826 407204
rect 317598 407192 317604 407204
rect 317656 407192 317662 407244
rect 151354 407124 151360 407176
rect 151412 407164 151418 407176
rect 161474 407164 161480 407176
rect 151412 407136 161480 407164
rect 151412 407124 151418 407136
rect 161474 407124 161480 407136
rect 161532 407124 161538 407176
rect 299382 407124 299388 407176
rect 299440 407164 299446 407176
rect 317506 407164 317512 407176
rect 299440 407136 317512 407164
rect 299440 407124 299446 407136
rect 317506 407124 317512 407136
rect 317564 407124 317570 407176
rect 52362 407056 52368 407108
rect 52420 407096 52426 407108
rect 166258 407096 166264 407108
rect 52420 407068 166264 407096
rect 52420 407056 52426 407068
rect 166258 407056 166264 407068
rect 166316 407056 166322 407108
rect 282822 407056 282828 407108
rect 282880 407096 282886 407108
rect 429470 407096 429476 407108
rect 282880 407068 429476 407096
rect 282880 407056 282886 407068
rect 429470 407056 429476 407068
rect 429528 407056 429534 407108
rect 56502 406988 56508 407040
rect 56560 407028 56566 407040
rect 170398 407028 170404 407040
rect 56560 407000 170404 407028
rect 56560 406988 56566 407000
rect 170398 406988 170404 407000
rect 170456 406988 170462 407040
rect 284110 406988 284116 407040
rect 284168 407028 284174 407040
rect 432690 407028 432696 407040
rect 284168 407000 432696 407028
rect 284168 406988 284174 407000
rect 432690 406988 432696 407000
rect 432748 406988 432754 407040
rect 59262 406920 59268 406972
rect 59320 406960 59326 406972
rect 173158 406960 173164 406972
rect 59320 406932 173164 406960
rect 59320 406920 59326 406932
rect 173158 406920 173164 406932
rect 173216 406920 173222 406972
rect 285582 406920 285588 406972
rect 285640 406960 285646 406972
rect 436186 406960 436192 406972
rect 285640 406932 436192 406960
rect 285640 406920 285646 406932
rect 436186 406920 436192 406932
rect 436244 406920 436250 406972
rect 53466 406852 53472 406904
rect 53524 406892 53530 406904
rect 169018 406892 169024 406904
rect 53524 406864 169024 406892
rect 53524 406852 53530 406864
rect 169018 406852 169024 406864
rect 169076 406852 169082 406904
rect 286962 406852 286968 406904
rect 287020 406892 287026 406904
rect 438946 406892 438952 406904
rect 287020 406864 438952 406892
rect 287020 406852 287026 406864
rect 438946 406852 438952 406864
rect 439004 406852 439010 406904
rect 61102 406784 61108 406836
rect 61160 406824 61166 406836
rect 178402 406824 178408 406836
rect 61160 406796 178408 406824
rect 61160 406784 61166 406796
rect 178402 406784 178408 406796
rect 178460 406784 178466 406836
rect 288342 406784 288348 406836
rect 288400 406824 288406 406836
rect 442166 406824 442172 406836
rect 288400 406796 442172 406824
rect 288400 406784 288406 406796
rect 442166 406784 442172 406796
rect 442224 406784 442230 406836
rect 99282 406716 99288 406768
rect 99340 406756 99346 406768
rect 332318 406756 332324 406768
rect 99340 406728 332324 406756
rect 99340 406716 99346 406728
rect 332318 406716 332324 406728
rect 332376 406716 332382 406768
rect 95970 406648 95976 406700
rect 96028 406688 96034 406700
rect 334986 406688 334992 406700
rect 96028 406660 334992 406688
rect 96028 406648 96034 406660
rect 334986 406648 334992 406660
rect 335044 406648 335050 406700
rect 86218 406580 86224 406632
rect 86276 406620 86282 406632
rect 326430 406620 326436 406632
rect 86276 406592 326436 406620
rect 86276 406580 86282 406592
rect 326430 406580 326436 406592
rect 326488 406580 326494 406632
rect 83642 406512 83648 406564
rect 83700 406552 83706 406564
rect 323946 406552 323952 406564
rect 83700 406524 323952 406552
rect 83700 406512 83706 406524
rect 323946 406512 323952 406524
rect 324004 406512 324010 406564
rect 88610 406444 88616 406496
rect 88668 406484 88674 406496
rect 336182 406484 336188 406496
rect 88668 406456 336188 406484
rect 88668 406444 88674 406456
rect 336182 406444 336188 406456
rect 336240 406444 336246 406496
rect 81066 406376 81072 406428
rect 81124 406416 81130 406428
rect 332134 406416 332140 406428
rect 81124 406388 332140 406416
rect 81124 406376 81130 406388
rect 332134 406376 332140 406388
rect 332192 406376 332198 406428
rect 48682 406308 48688 406360
rect 48740 406348 48746 406360
rect 162118 406348 162124 406360
rect 48740 406320 162124 406348
rect 48740 406308 48746 406320
rect 162118 406308 162124 406320
rect 162176 406308 162182 406360
rect 281442 406308 281448 406360
rect 281500 406348 281506 406360
rect 426434 406348 426440 406360
rect 281500 406320 426440 406348
rect 281500 406308 281506 406320
rect 426434 406308 426440 406320
rect 426492 406308 426498 406360
rect 278590 406240 278596 406292
rect 278648 406280 278654 406292
rect 423766 406280 423772 406292
rect 278648 406252 423772 406280
rect 278648 406240 278654 406252
rect 423766 406240 423772 406252
rect 423824 406240 423830 406292
rect 277302 406172 277308 406224
rect 277360 406212 277366 406224
rect 419994 406212 420000 406224
rect 277360 406184 420000 406212
rect 277360 406172 277366 406184
rect 419994 406172 420000 406184
rect 420052 406172 420058 406224
rect 275922 406104 275928 406156
rect 275980 406144 275986 406156
rect 416866 406144 416872 406156
rect 275980 406116 416872 406144
rect 275980 406104 275986 406116
rect 416866 406104 416872 406116
rect 416924 406104 416930 406156
rect 242802 406036 242808 406088
rect 242860 406076 242866 406088
rect 353662 406076 353668 406088
rect 242860 406048 353668 406076
rect 242860 406036 242866 406048
rect 353662 406036 353668 406048
rect 353720 406036 353726 406088
rect 241330 405968 241336 406020
rect 241388 406008 241394 406020
rect 349430 406008 349436 406020
rect 241388 405980 349436 406008
rect 241388 405968 241394 405980
rect 349430 405968 349436 405980
rect 349488 405968 349494 406020
rect 238570 405900 238576 405952
rect 238628 405940 238634 405952
rect 322382 405940 322388 405952
rect 238628 405912 322388 405940
rect 238628 405900 238634 405912
rect 322382 405900 322388 405912
rect 322440 405900 322446 405952
rect 243722 405832 243728 405884
rect 243780 405872 243786 405884
rect 321278 405872 321284 405884
rect 243780 405844 321284 405872
rect 243780 405832 243786 405844
rect 321278 405832 321284 405844
rect 321336 405832 321342 405884
rect 281074 405764 281080 405816
rect 281132 405804 281138 405816
rect 318334 405804 318340 405816
rect 281132 405776 318340 405804
rect 281132 405764 281138 405776
rect 318334 405764 318340 405776
rect 318392 405764 318398 405816
rect 397362 403656 397368 403708
rect 397420 403696 397426 403708
rect 503714 403696 503720 403708
rect 397420 403668 503720 403696
rect 397420 403656 397426 403668
rect 503714 403656 503720 403668
rect 503772 403656 503778 403708
rect 394418 403588 394424 403640
rect 394476 403628 394482 403640
rect 502334 403628 502340 403640
rect 394476 403600 502340 403628
rect 394476 403588 394482 403600
rect 502334 403588 502340 403600
rect 502392 403588 502398 403640
rect 400766 402500 400772 402552
rect 400824 402540 400830 402552
rect 506474 402540 506480 402552
rect 400824 402512 506480 402540
rect 400824 402500 400830 402512
rect 506474 402500 506480 402512
rect 506532 402500 506538 402552
rect 391290 402432 391296 402484
rect 391348 402472 391354 402484
rect 500954 402472 500960 402484
rect 391348 402444 500960 402472
rect 391348 402432 391354 402444
rect 500954 402432 500960 402444
rect 501012 402432 501018 402484
rect 388070 402364 388076 402416
rect 388128 402404 388134 402416
rect 499574 402404 499580 402416
rect 388128 402376 499580 402404
rect 388128 402364 388134 402376
rect 499574 402364 499580 402376
rect 499632 402364 499638 402416
rect 384942 402296 384948 402348
rect 385000 402336 385006 402348
rect 497458 402336 497464 402348
rect 385000 402308 497464 402336
rect 385000 402296 385006 402308
rect 497458 402296 497464 402308
rect 497516 402296 497522 402348
rect 375282 402228 375288 402280
rect 375340 402268 375346 402280
rect 492674 402268 492680 402280
rect 375340 402240 492680 402268
rect 375340 402228 375346 402240
rect 492674 402228 492680 402240
rect 492732 402228 492738 402280
rect 320082 401616 320088 401668
rect 320140 401656 320146 401668
rect 323762 401656 323768 401668
rect 320140 401628 323768 401656
rect 320140 401616 320146 401628
rect 323762 401616 323768 401628
rect 323820 401616 323826 401668
rect 349062 401548 349068 401600
rect 349120 401588 349126 401600
rect 420178 401588 420184 401600
rect 349120 401560 420184 401588
rect 349120 401548 349126 401560
rect 420178 401548 420184 401560
rect 420236 401548 420242 401600
rect 421558 401548 421564 401600
rect 421616 401588 421622 401600
rect 433794 401588 433800 401600
rect 421616 401560 433800 401588
rect 421616 401548 421622 401560
rect 433794 401548 433800 401560
rect 433852 401548 433858 401600
rect 443638 401588 443644 401600
rect 441586 401560 443644 401588
rect 341518 401480 341524 401532
rect 341576 401520 341582 401532
rect 347866 401520 347872 401532
rect 341576 401492 347872 401520
rect 341576 401480 341582 401492
rect 347866 401480 347872 401492
rect 347924 401480 347930 401532
rect 353202 401480 353208 401532
rect 353260 401520 353266 401532
rect 441586 401520 441614 401560
rect 443638 401548 443644 401560
rect 443696 401548 443702 401600
rect 451090 401548 451096 401600
rect 451148 401588 451154 401600
rect 472250 401588 472256 401600
rect 451148 401560 472256 401588
rect 451148 401548 451154 401560
rect 472250 401548 472256 401560
rect 472308 401548 472314 401600
rect 353260 401492 441614 401520
rect 353260 401480 353266 401492
rect 449158 401480 449164 401532
rect 449216 401520 449222 401532
rect 465905 401523 465963 401529
rect 449216 401492 465856 401520
rect 449216 401480 449222 401492
rect 334710 401412 334716 401464
rect 334768 401452 334774 401464
rect 370590 401452 370596 401464
rect 334768 401424 370596 401452
rect 334768 401412 334774 401424
rect 370590 401412 370596 401424
rect 370648 401412 370654 401464
rect 378781 401455 378839 401461
rect 378781 401421 378793 401455
rect 378827 401452 378839 401455
rect 465721 401455 465779 401461
rect 465721 401452 465733 401455
rect 378827 401424 465733 401452
rect 378827 401421 378839 401424
rect 378781 401415 378839 401421
rect 465721 401421 465733 401424
rect 465767 401421 465779 401455
rect 465721 401415 465779 401421
rect 323578 401344 323584 401396
rect 323636 401384 323642 401396
rect 440234 401384 440240 401396
rect 323636 401356 440240 401384
rect 323636 401344 323642 401356
rect 440234 401344 440240 401356
rect 440292 401344 440298 401396
rect 447042 401344 447048 401396
rect 447100 401384 447106 401396
rect 465828 401384 465856 401492
rect 465905 401489 465917 401523
rect 465951 401520 465963 401523
rect 465951 401492 470594 401520
rect 465951 401489 465963 401492
rect 465905 401483 465963 401489
rect 470566 401452 470594 401492
rect 482278 401452 482284 401464
rect 470566 401424 482284 401452
rect 482278 401412 482284 401424
rect 482336 401412 482342 401464
rect 472342 401384 472348 401396
rect 447100 401356 465764 401384
rect 465828 401356 472348 401384
rect 447100 401344 447106 401356
rect 324958 401276 324964 401328
rect 325016 401316 325022 401328
rect 443270 401316 443276 401328
rect 325016 401288 443276 401316
rect 325016 401276 325022 401288
rect 443270 401276 443276 401288
rect 443328 401276 443334 401328
rect 446030 401276 446036 401328
rect 446088 401316 446094 401328
rect 465629 401319 465687 401325
rect 465629 401316 465641 401319
rect 446088 401288 465641 401316
rect 446088 401276 446094 401288
rect 465629 401285 465641 401288
rect 465675 401285 465687 401319
rect 465736 401316 465764 401356
rect 472342 401344 472348 401356
rect 472400 401344 472406 401396
rect 472526 401316 472532 401328
rect 465736 401288 472532 401316
rect 465629 401279 465687 401285
rect 472526 401276 472532 401288
rect 472584 401276 472590 401328
rect 342898 401208 342904 401260
rect 342956 401248 342962 401260
rect 346394 401248 346400 401260
rect 342956 401220 346400 401248
rect 342956 401208 342962 401220
rect 346394 401208 346400 401220
rect 346452 401208 346458 401260
rect 353938 401208 353944 401260
rect 353996 401248 354002 401260
rect 360194 401248 360200 401260
rect 353996 401220 360200 401248
rect 353996 401208 354002 401220
rect 360194 401208 360200 401220
rect 360252 401208 360258 401260
rect 362862 401208 362868 401260
rect 362920 401248 362926 401260
rect 480898 401248 480904 401260
rect 362920 401220 480904 401248
rect 362920 401208 362926 401220
rect 480898 401208 480904 401220
rect 480956 401208 480962 401260
rect 327718 401140 327724 401192
rect 327776 401180 327782 401192
rect 354950 401180 354956 401192
rect 327776 401152 354956 401180
rect 327776 401140 327782 401152
rect 354950 401140 354956 401152
rect 355008 401140 355014 401192
rect 369121 401183 369179 401189
rect 369121 401149 369133 401183
rect 369167 401180 369179 401183
rect 478138 401180 478144 401192
rect 369167 401152 478144 401180
rect 369167 401149 369179 401152
rect 369121 401143 369179 401149
rect 478138 401140 478144 401152
rect 478196 401140 478202 401192
rect 322198 401072 322204 401124
rect 322256 401112 322262 401124
rect 350626 401112 350632 401124
rect 322256 401084 350632 401112
rect 322256 401072 322262 401084
rect 350626 401072 350632 401084
rect 350684 401072 350690 401124
rect 356514 401072 356520 401124
rect 356572 401112 356578 401124
rect 476758 401112 476764 401124
rect 356572 401084 476764 401112
rect 356572 401072 356578 401084
rect 476758 401072 476764 401084
rect 476816 401072 476822 401124
rect 343910 401004 343916 401056
rect 343968 401044 343974 401056
rect 474734 401044 474740 401056
rect 343968 401016 474740 401044
rect 343968 401004 343974 401016
rect 474734 401004 474740 401016
rect 474792 401004 474798 401056
rect 316678 400936 316684 400988
rect 316736 400976 316742 400988
rect 455874 400976 455880 400988
rect 316736 400948 455880 400976
rect 316736 400936 316742 400948
rect 455874 400936 455880 400948
rect 455932 400936 455938 400988
rect 465629 400979 465687 400985
rect 465629 400945 465641 400979
rect 465675 400976 465687 400979
rect 472434 400976 472440 400988
rect 465675 400948 472440 400976
rect 465675 400945 465687 400948
rect 465629 400939 465687 400945
rect 472434 400936 472440 400948
rect 472492 400936 472498 400988
rect 316770 400868 316776 400920
rect 316828 400908 316834 400920
rect 456978 400908 456984 400920
rect 316828 400880 456984 400908
rect 316828 400868 316834 400880
rect 456978 400868 456984 400880
rect 457036 400868 457042 400920
rect 478690 400868 478696 400920
rect 478748 400908 478754 400920
rect 530578 400908 530584 400920
rect 478748 400880 530584 400908
rect 478748 400868 478754 400880
rect 530578 400868 530584 400880
rect 530636 400868 530642 400920
rect 344738 400800 344744 400852
rect 344796 400840 344802 400852
rect 409138 400840 409144 400852
rect 344796 400812 409144 400840
rect 344796 400800 344802 400812
rect 409138 400800 409144 400812
rect 409196 400800 409202 400852
rect 410610 400800 410616 400852
rect 410668 400840 410674 400852
rect 427814 400840 427820 400852
rect 410668 400812 427820 400840
rect 410668 400800 410674 400812
rect 427814 400800 427820 400812
rect 427872 400800 427878 400852
rect 431218 400800 431224 400852
rect 431276 400840 431282 400852
rect 436922 400840 436928 400852
rect 431276 400812 436928 400840
rect 431276 400800 431282 400812
rect 436922 400800 436928 400812
rect 436980 400800 436986 400852
rect 453390 400800 453396 400852
rect 453448 400840 453454 400852
rect 472158 400840 472164 400852
rect 453448 400812 472164 400840
rect 453448 400800 453454 400812
rect 472158 400800 472164 400812
rect 472216 400800 472222 400852
rect 349798 400732 349804 400784
rect 349856 400772 349862 400784
rect 363230 400772 363236 400784
rect 349856 400744 363236 400772
rect 349856 400732 349862 400744
rect 363230 400732 363236 400744
rect 363288 400732 363294 400784
rect 363598 400732 363604 400784
rect 363656 400772 363662 400784
rect 418154 400772 418160 400784
rect 363656 400744 418160 400772
rect 363656 400732 363662 400744
rect 418154 400732 418160 400744
rect 418212 400732 418218 400784
rect 331950 400664 331956 400716
rect 332008 400704 332014 400716
rect 364518 400704 364524 400716
rect 332008 400676 364524 400704
rect 332008 400664 332014 400676
rect 364518 400664 364524 400676
rect 364576 400664 364582 400716
rect 372338 400664 372344 400716
rect 372396 400704 372402 400716
rect 378781 400707 378839 400713
rect 378781 400704 378793 400707
rect 372396 400676 378793 400704
rect 372396 400664 372402 400676
rect 378781 400673 378793 400676
rect 378827 400673 378839 400707
rect 378781 400667 378839 400673
rect 382918 400664 382924 400716
rect 382976 400704 382982 400716
rect 408494 400704 408500 400716
rect 382976 400676 408500 400704
rect 382976 400664 382982 400676
rect 408494 400664 408500 400676
rect 408552 400664 408558 400716
rect 417418 400664 417424 400716
rect 417476 400704 417482 400716
rect 430666 400704 430672 400716
rect 417476 400676 430672 400704
rect 417476 400664 417482 400676
rect 430666 400664 430672 400676
rect 430724 400664 430730 400716
rect 359642 400596 359648 400648
rect 359700 400636 359706 400648
rect 369121 400639 369179 400645
rect 369121 400636 369133 400639
rect 359700 400608 369133 400636
rect 359700 400596 359706 400608
rect 369121 400605 369133 400608
rect 369167 400605 369179 400639
rect 369121 400599 369179 400605
rect 370498 400596 370504 400648
rect 370556 400636 370562 400648
rect 382274 400636 382280 400648
rect 370556 400608 382280 400636
rect 370556 400596 370562 400608
rect 382274 400596 382280 400608
rect 382332 400596 382338 400648
rect 395338 400596 395344 400648
rect 395396 400636 395402 400648
rect 414842 400636 414848 400648
rect 395396 400608 414848 400636
rect 395396 400596 395402 400608
rect 414842 400596 414848 400608
rect 414900 400596 414906 400648
rect 399478 400460 399484 400512
rect 399536 400500 399542 400512
rect 411714 400500 411720 400512
rect 399536 400472 411720 400500
rect 399536 400460 399542 400472
rect 411714 400460 411720 400472
rect 411772 400460 411778 400512
rect 413278 400460 413284 400512
rect 413336 400500 413342 400512
rect 424318 400500 424324 400512
rect 413336 400472 424324 400500
rect 413336 400460 413342 400472
rect 424318 400460 424324 400472
rect 424376 400460 424382 400512
rect 407758 400324 407764 400376
rect 407816 400364 407822 400376
rect 421190 400364 421196 400376
rect 407816 400336 421196 400364
rect 407816 400324 407822 400336
rect 421190 400324 421196 400336
rect 421248 400324 421254 400376
rect 472802 400324 472808 400376
rect 472860 400364 472866 400376
rect 476942 400364 476948 400376
rect 472860 400336 476948 400364
rect 472860 400324 472866 400336
rect 476942 400324 476948 400336
rect 477000 400324 477006 400376
rect 364978 400256 364984 400308
rect 365036 400296 365042 400308
rect 366450 400296 366456 400308
rect 365036 400268 366456 400296
rect 365036 400256 365042 400268
rect 366450 400256 366456 400268
rect 366508 400256 366514 400308
rect 393958 400256 393964 400308
rect 394016 400296 394022 400308
rect 402238 400296 402244 400308
rect 394016 400268 402244 400296
rect 394016 400256 394022 400268
rect 402238 400256 402244 400268
rect 402296 400256 402302 400308
rect 472710 400256 472716 400308
rect 472768 400296 472774 400308
rect 474826 400296 474832 400308
rect 472768 400268 474832 400296
rect 472768 400256 472774 400268
rect 474826 400256 474832 400268
rect 474884 400256 474890 400308
rect 365990 400188 365996 400240
rect 366048 400228 366054 400240
rect 367002 400228 367008 400240
rect 366048 400200 367008 400228
rect 366048 400188 366054 400200
rect 367002 400188 367008 400200
rect 367060 400188 367066 400240
rect 369118 400188 369124 400240
rect 369176 400228 369182 400240
rect 369762 400228 369768 400240
rect 369176 400200 369768 400228
rect 369176 400188 369182 400200
rect 369762 400188 369768 400200
rect 369820 400188 369826 400240
rect 371878 400188 371884 400240
rect 371936 400228 371942 400240
rect 372706 400228 372712 400240
rect 371936 400200 372712 400228
rect 371936 400188 371942 400200
rect 372706 400188 372712 400200
rect 372764 400188 372770 400240
rect 374638 400188 374644 400240
rect 374696 400228 374702 400240
rect 375926 400228 375932 400240
rect 374696 400200 375932 400228
rect 374696 400188 374702 400200
rect 375926 400188 375932 400200
rect 375984 400188 375990 400240
rect 378594 400188 378600 400240
rect 378652 400228 378658 400240
rect 379422 400228 379428 400240
rect 378652 400200 379428 400228
rect 378652 400188 378658 400200
rect 379422 400188 379428 400200
rect 379480 400188 379486 400240
rect 388438 400188 388444 400240
rect 388496 400228 388502 400240
rect 392026 400228 392032 400240
rect 388496 400200 392032 400228
rect 388496 400188 388502 400200
rect 392026 400188 392032 400200
rect 392084 400188 392090 400240
rect 396718 400188 396724 400240
rect 396776 400228 396782 400240
rect 398006 400228 398012 400240
rect 396776 400200 398012 400228
rect 396776 400188 396782 400200
rect 398006 400188 398012 400200
rect 398064 400188 398070 400240
rect 403618 400188 403624 400240
rect 403676 400228 403682 400240
rect 404354 400228 404360 400240
rect 403676 400200 404360 400228
rect 403676 400188 403682 400200
rect 404354 400188 404360 400200
rect 404412 400188 404418 400240
rect 410242 400188 410248 400240
rect 410300 400228 410306 400240
rect 411898 400228 411904 400240
rect 410300 400200 411904 400228
rect 410300 400188 410306 400200
rect 411898 400188 411904 400200
rect 411956 400188 411962 400240
rect 413370 400188 413376 400240
rect 413428 400228 413434 400240
rect 414658 400228 414664 400240
rect 413428 400200 414664 400228
rect 413428 400188 413434 400200
rect 414658 400188 414664 400200
rect 414716 400188 414722 400240
rect 422846 400188 422852 400240
rect 422904 400228 422910 400240
rect 423582 400228 423588 400240
rect 422904 400200 423588 400228
rect 422904 400188 422910 400200
rect 423582 400188 423588 400200
rect 423640 400188 423646 400240
rect 432322 400188 432328 400240
rect 432380 400228 432386 400240
rect 433242 400228 433248 400240
rect 432380 400200 433248 400228
rect 432380 400188 432386 400200
rect 433242 400188 433248 400200
rect 433300 400188 433306 400240
rect 435450 400188 435456 400240
rect 435508 400228 435514 400240
rect 436002 400228 436008 400240
rect 435508 400200 436008 400228
rect 435508 400188 435514 400200
rect 436002 400188 436008 400200
rect 436060 400188 436066 400240
rect 458634 400188 458640 400240
rect 458692 400228 458698 400240
rect 459462 400228 459468 400240
rect 458692 400200 459468 400228
rect 458692 400188 458698 400200
rect 459462 400188 459468 400200
rect 459520 400188 459526 400240
rect 472894 400188 472900 400240
rect 472952 400228 472958 400240
rect 473814 400228 473820 400240
rect 472952 400200 473820 400228
rect 472952 400188 472958 400200
rect 473814 400188 473820 400200
rect 473872 400188 473878 400240
rect 475378 400188 475384 400240
rect 475436 400228 475442 400240
rect 476114 400228 476120 400240
rect 475436 400200 476120 400228
rect 475436 400188 475442 400200
rect 476114 400188 476120 400200
rect 476172 400188 476178 400240
rect 479702 400188 479708 400240
rect 479760 400228 479766 400240
rect 480162 400228 480168 400240
rect 479760 400200 480168 400228
rect 479760 400188 479766 400200
rect 480162 400188 480168 400200
rect 480220 400188 480226 400240
rect 462314 400120 462320 400172
rect 462372 400160 462378 400172
rect 463234 400160 463240 400172
rect 462372 400132 463240 400160
rect 462372 400120 462378 400132
rect 463234 400120 463240 400132
rect 463292 400120 463298 400172
rect 467834 400120 467840 400172
rect 467892 400160 467898 400172
rect 468570 400160 468576 400172
rect 467892 400132 468576 400160
rect 467892 400120 467898 400132
rect 468570 400120 468576 400132
rect 468628 400120 468634 400172
rect 320818 397468 320824 397520
rect 320876 397508 320882 397520
rect 337654 397508 337660 397520
rect 320876 397480 337660 397508
rect 320876 397468 320882 397480
rect 337654 397468 337660 397480
rect 337712 397468 337718 397520
rect 322198 396040 322204 396092
rect 322256 396080 322262 396092
rect 337654 396080 337660 396092
rect 322256 396052 337660 396080
rect 322256 396040 322262 396052
rect 337654 396040 337660 396052
rect 337712 396040 337718 396092
rect 482922 395972 482928 396024
rect 482980 396012 482986 396024
rect 536098 396012 536104 396024
rect 482980 395984 536104 396012
rect 482980 395972 482986 395984
rect 536098 395972 536104 395984
rect 536156 395972 536162 396024
rect 329098 394748 329104 394800
rect 329156 394788 329162 394800
rect 337654 394788 337660 394800
rect 329156 394760 337660 394788
rect 329156 394748 329162 394760
rect 337654 394748 337660 394760
rect 337712 394748 337718 394800
rect 321186 394680 321192 394732
rect 321244 394720 321250 394732
rect 337746 394720 337752 394732
rect 321244 394692 337752 394720
rect 321244 394680 321250 394692
rect 337746 394680 337752 394692
rect 337804 394680 337810 394732
rect 330478 393388 330484 393440
rect 330536 393428 330542 393440
rect 337654 393428 337660 393440
rect 330536 393400 337660 393428
rect 330536 393388 330542 393400
rect 337654 393388 337660 393400
rect 337712 393388 337718 393440
rect 323578 393320 323584 393372
rect 323636 393360 323642 393372
rect 337746 393360 337752 393372
rect 323636 393332 337752 393360
rect 323636 393320 323642 393332
rect 337746 393320 337752 393332
rect 337804 393320 337810 393372
rect 331950 392028 331956 392080
rect 332008 392068 332014 392080
rect 337654 392068 337660 392080
rect 332008 392040 337660 392068
rect 332008 392028 332014 392040
rect 337654 392028 337660 392040
rect 337712 392028 337718 392080
rect 325050 391960 325056 392012
rect 325108 392000 325114 392012
rect 337746 392000 337752 392012
rect 325108 391972 337752 392000
rect 325108 391960 325114 391972
rect 337746 391960 337752 391972
rect 337804 391960 337810 392012
rect 482922 391892 482928 391944
rect 482980 391932 482986 391944
rect 529198 391932 529204 391944
rect 482980 391904 529204 391932
rect 482980 391892 482986 391904
rect 529198 391892 529204 391904
rect 529256 391892 529262 391944
rect 334710 390600 334716 390652
rect 334768 390640 334774 390652
rect 337654 390640 337660 390652
rect 334768 390612 337660 390640
rect 334768 390600 334774 390612
rect 337654 390600 337660 390612
rect 337712 390600 337718 390652
rect 324958 390532 324964 390584
rect 325016 390572 325022 390584
rect 337746 390572 337752 390584
rect 325016 390544 337752 390572
rect 325016 390532 325022 390544
rect 337746 390532 337752 390544
rect 337804 390532 337810 390584
rect 328086 389308 328092 389360
rect 328144 389348 328150 389360
rect 337654 389348 337660 389360
rect 328144 389320 337660 389348
rect 328144 389308 328150 389320
rect 337654 389308 337660 389320
rect 337712 389308 337718 389360
rect 327718 389240 327724 389292
rect 327776 389280 327782 389292
rect 337746 389280 337752 389292
rect 327776 389252 337752 389280
rect 327776 389240 327782 389252
rect 337746 389240 337752 389252
rect 337804 389240 337810 389292
rect 322474 389172 322480 389224
rect 322532 389212 322538 389224
rect 337654 389212 337660 389224
rect 322532 389184 337660 389212
rect 322532 389172 322538 389184
rect 337654 389172 337660 389184
rect 337712 389172 337718 389224
rect 316862 389104 316868 389156
rect 316920 389144 316926 389156
rect 337838 389144 337844 389156
rect 316920 389116 337844 389144
rect 316920 389104 316926 389116
rect 337838 389104 337844 389116
rect 337896 389104 337902 389156
rect 318150 389036 318156 389088
rect 318208 389076 318214 389088
rect 337746 389076 337752 389088
rect 318208 389048 337752 389076
rect 318208 389036 318214 389048
rect 337746 389036 337752 389048
rect 337804 389036 337810 389088
rect 328270 387744 328276 387796
rect 328328 387784 328334 387796
rect 337654 387784 337660 387796
rect 328328 387756 337660 387784
rect 328328 387744 328334 387756
rect 337654 387744 337660 387756
rect 337712 387744 337718 387796
rect 329558 387676 329564 387728
rect 329616 387716 329622 387728
rect 337746 387716 337752 387728
rect 329616 387688 337752 387716
rect 329616 387676 329622 387688
rect 337746 387676 337752 387688
rect 337804 387676 337810 387728
rect 325326 386316 325332 386368
rect 325384 386356 325390 386368
rect 337654 386356 337660 386368
rect 325384 386328 337660 386356
rect 325384 386316 325390 386328
rect 337654 386316 337660 386328
rect 337712 386316 337718 386368
rect 482922 386316 482928 386368
rect 482980 386356 482986 386368
rect 533338 386356 533344 386368
rect 482980 386328 533344 386356
rect 482980 386316 482986 386328
rect 533338 386316 533344 386328
rect 533396 386316 533402 386368
rect 330570 386044 330576 386096
rect 330628 386084 330634 386096
rect 337746 386084 337752 386096
rect 330628 386056 337752 386084
rect 330628 386044 330634 386056
rect 337746 386044 337752 386056
rect 337804 386044 337810 386096
rect 320910 384956 320916 385008
rect 320968 384996 320974 385008
rect 337654 384996 337660 385008
rect 320968 384968 337660 384996
rect 320968 384956 320974 384968
rect 337654 384956 337660 384968
rect 337712 384956 337718 385008
rect 322750 384888 322756 384940
rect 322808 384928 322814 384940
rect 337746 384928 337752 384940
rect 322808 384900 337752 384928
rect 322808 384888 322814 384900
rect 337746 384888 337752 384900
rect 337804 384888 337810 384940
rect 322290 383596 322296 383648
rect 322348 383636 322354 383648
rect 337654 383636 337660 383648
rect 322348 383608 337660 383636
rect 322348 383596 322354 383608
rect 337654 383596 337660 383608
rect 337712 383596 337718 383648
rect 334618 383528 334624 383580
rect 334676 383568 334682 383580
rect 337746 383568 337752 383580
rect 334676 383540 337752 383568
rect 334676 383528 334682 383540
rect 337746 383528 337752 383540
rect 337804 383528 337810 383580
rect 331858 382168 331864 382220
rect 331916 382208 331922 382220
rect 336918 382208 336924 382220
rect 331916 382180 336924 382208
rect 331916 382168 331922 382180
rect 336918 382168 336924 382180
rect 336976 382168 336982 382220
rect 482002 382168 482008 382220
rect 482060 382208 482066 382220
rect 538858 382208 538864 382220
rect 482060 382180 538864 382208
rect 482060 382168 482066 382180
rect 538858 382168 538864 382180
rect 538916 382168 538922 382220
rect 330938 382100 330944 382152
rect 330996 382140 331002 382152
rect 337654 382140 337660 382152
rect 330996 382112 337660 382140
rect 330996 382100 331002 382112
rect 337654 382100 337660 382112
rect 337712 382100 337718 382152
rect 323670 380740 323676 380792
rect 323728 380780 323734 380792
rect 337746 380780 337752 380792
rect 323728 380752 337752 380780
rect 323728 380740 323734 380752
rect 337746 380740 337752 380752
rect 337804 380740 337810 380792
rect 319438 380672 319444 380724
rect 319496 380712 319502 380724
rect 336918 380712 336924 380724
rect 319496 380684 336924 380712
rect 319496 380672 319502 380684
rect 336918 380672 336924 380684
rect 336976 380672 336982 380724
rect 329466 379448 329472 379500
rect 329524 379488 329530 379500
rect 337746 379488 337752 379500
rect 329524 379460 337752 379488
rect 329524 379448 329530 379460
rect 337746 379448 337752 379460
rect 337804 379448 337810 379500
rect 319438 378156 319444 378208
rect 319496 378196 319502 378208
rect 337654 378196 337660 378208
rect 319496 378168 337660 378196
rect 319496 378156 319502 378168
rect 337654 378156 337660 378168
rect 337712 378156 337718 378208
rect 482186 378156 482192 378208
rect 482244 378196 482250 378208
rect 580166 378196 580172 378208
rect 482244 378168 580172 378196
rect 482244 378156 482250 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 327994 378088 328000 378140
rect 328052 378128 328058 378140
rect 337746 378128 337752 378140
rect 328052 378100 337752 378128
rect 328052 378088 328058 378100
rect 337746 378088 337752 378100
rect 337804 378088 337810 378140
rect 482278 378088 482284 378140
rect 482336 378128 482342 378140
rect 580258 378128 580264 378140
rect 482336 378100 580264 378128
rect 482336 378088 482342 378100
rect 580258 378088 580264 378100
rect 580316 378088 580322 378140
rect 318150 376728 318156 376780
rect 318208 376768 318214 376780
rect 337286 376768 337292 376780
rect 318208 376740 337292 376768
rect 318208 376728 318214 376740
rect 337286 376728 337292 376740
rect 337344 376728 337350 376780
rect 318242 376660 318248 376712
rect 318300 376700 318306 376712
rect 337654 376700 337660 376712
rect 318300 376672 337660 376700
rect 318300 376660 318306 376672
rect 337654 376660 337660 376672
rect 337712 376660 337718 376712
rect 330570 375368 330576 375420
rect 330628 375408 330634 375420
rect 337102 375408 337108 375420
rect 330628 375380 337108 375408
rect 330628 375368 330634 375380
rect 337102 375368 337108 375380
rect 337160 375368 337166 375420
rect 318334 375300 318340 375352
rect 318392 375340 318398 375352
rect 337654 375340 337660 375352
rect 318392 375312 337660 375340
rect 318392 375300 318398 375312
rect 337654 375300 337660 375312
rect 337712 375300 337718 375352
rect 318242 374008 318248 374060
rect 318300 374048 318306 374060
rect 337746 374048 337752 374060
rect 318300 374020 337752 374048
rect 318300 374008 318306 374020
rect 337746 374008 337752 374020
rect 337804 374008 337810 374060
rect 322658 373940 322664 373992
rect 322716 373980 322722 373992
rect 337654 373980 337660 373992
rect 322716 373952 337660 373980
rect 322716 373940 322722 373952
rect 337654 373940 337660 373952
rect 337712 373940 337718 373992
rect 326614 372580 326620 372632
rect 326672 372620 326678 372632
rect 337746 372620 337752 372632
rect 326672 372592 337752 372620
rect 326672 372580 326678 372592
rect 337746 372580 337752 372592
rect 337804 372580 337810 372632
rect 482922 372512 482928 372564
rect 482980 372552 482986 372564
rect 537478 372552 537484 372564
rect 482980 372524 537484 372552
rect 482980 372512 482986 372524
rect 537478 372512 537484 372524
rect 537536 372512 537542 372564
rect 318426 371832 318432 371884
rect 318484 371872 318490 371884
rect 318484 371844 335354 371872
rect 318484 371832 318490 371844
rect 335326 371804 335354 371844
rect 337562 371804 337568 371816
rect 335326 371776 337568 371804
rect 337562 371764 337568 371776
rect 337620 371764 337626 371816
rect 318334 371220 318340 371272
rect 318392 371260 318398 371272
rect 336918 371260 336924 371272
rect 318392 371232 336924 371260
rect 318392 371220 318398 371232
rect 336918 371220 336924 371232
rect 336976 371220 336982 371272
rect 321370 371152 321376 371204
rect 321428 371192 321434 371204
rect 337654 371192 337660 371204
rect 321428 371164 337660 371192
rect 321428 371152 321434 371164
rect 337654 371152 337660 371164
rect 337712 371152 337718 371204
rect 318426 369860 318432 369912
rect 318484 369900 318490 369912
rect 337654 369900 337660 369912
rect 318484 369872 337660 369900
rect 318484 369860 318490 369872
rect 337654 369860 337660 369872
rect 337712 369860 337718 369912
rect 322566 369792 322572 369844
rect 322624 369832 322630 369844
rect 337286 369832 337292 369844
rect 322624 369804 337292 369832
rect 322624 369792 322630 369804
rect 337286 369792 337292 369804
rect 337344 369792 337350 369844
rect 333422 368500 333428 368552
rect 333480 368540 333486 368552
rect 337654 368540 337660 368552
rect 333480 368512 337660 368540
rect 333480 368500 333486 368512
rect 337654 368500 337660 368512
rect 337712 368500 337718 368552
rect 318518 368432 318524 368484
rect 318576 368472 318582 368484
rect 337746 368472 337752 368484
rect 318576 368444 337752 368472
rect 318576 368432 318582 368444
rect 337746 368432 337752 368444
rect 337804 368432 337810 368484
rect 329466 367072 329472 367124
rect 329524 367112 329530 367124
rect 337746 367112 337752 367124
rect 329524 367084 337752 367112
rect 329524 367072 329530 367084
rect 337746 367072 337752 367084
rect 337804 367072 337810 367124
rect 335170 365712 335176 365764
rect 335228 365752 335234 365764
rect 337286 365752 337292 365764
rect 335228 365724 337292 365752
rect 335228 365712 335234 365724
rect 337286 365712 337292 365724
rect 337344 365712 337350 365764
rect 332410 365644 332416 365696
rect 332468 365684 332474 365696
rect 337654 365684 337660 365696
rect 332468 365656 337660 365684
rect 332468 365644 332474 365656
rect 337654 365644 337660 365656
rect 337712 365644 337718 365696
rect 327994 364352 328000 364404
rect 328052 364392 328058 364404
rect 337746 364392 337752 364404
rect 328052 364364 337752 364392
rect 328052 364352 328058 364364
rect 337746 364352 337752 364364
rect 337804 364352 337810 364404
rect 482370 364352 482376 364404
rect 482428 364392 482434 364404
rect 580166 364392 580172 364404
rect 482428 364364 580172 364392
rect 482428 364352 482434 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 335262 364284 335268 364336
rect 335320 364324 335326 364336
rect 337654 364324 337660 364336
rect 335320 364296 337660 364324
rect 335320 364284 335326 364296
rect 337654 364284 337660 364296
rect 337712 364284 337718 364336
rect 322566 362924 322572 362976
rect 322624 362964 322630 362976
rect 337746 362964 337752 362976
rect 322624 362936 337752 362964
rect 322624 362924 322630 362936
rect 337746 362924 337752 362936
rect 337804 362924 337810 362976
rect 328178 362856 328184 362908
rect 328236 362896 328242 362908
rect 337654 362896 337660 362908
rect 328236 362868 337660 362896
rect 328236 362856 328242 362868
rect 337654 362856 337660 362868
rect 337712 362856 337718 362908
rect 322290 361564 322296 361616
rect 322348 361604 322354 361616
rect 337102 361604 337108 361616
rect 322348 361576 337108 361604
rect 322348 361564 322354 361576
rect 337102 361564 337108 361576
rect 337160 361564 337166 361616
rect 325510 361496 325516 361548
rect 325568 361536 325574 361548
rect 336918 361536 336924 361548
rect 325568 361508 336924 361536
rect 325568 361496 325574 361508
rect 336918 361496 336924 361508
rect 336976 361496 336982 361548
rect 329558 360204 329564 360256
rect 329616 360244 329622 360256
rect 337654 360244 337660 360256
rect 329616 360216 337660 360244
rect 329616 360204 329622 360216
rect 337654 360204 337660 360216
rect 337712 360204 337718 360256
rect 319622 359456 319628 359508
rect 319680 359496 319686 359508
rect 337562 359496 337568 359508
rect 319680 359468 337568 359496
rect 319680 359456 319686 359468
rect 337562 359456 337568 359468
rect 337620 359456 337626 359508
rect 320910 358776 320916 358828
rect 320968 358816 320974 358828
rect 337654 358816 337660 358828
rect 320968 358788 337660 358816
rect 320968 358776 320974 358788
rect 337654 358776 337660 358788
rect 337712 358776 337718 358828
rect 335078 358708 335084 358760
rect 335136 358748 335142 358760
rect 336918 358748 336924 358760
rect 335136 358720 336924 358748
rect 335136 358708 335142 358720
rect 336918 358708 336924 358720
rect 336976 358708 336982 358760
rect 325326 357416 325332 357468
rect 325384 357456 325390 357468
rect 337746 357456 337752 357468
rect 325384 357428 337752 357456
rect 325384 357416 325390 357428
rect 337746 357416 337752 357428
rect 337804 357416 337810 357468
rect 319530 357348 319536 357400
rect 319588 357388 319594 357400
rect 337654 357388 337660 357400
rect 319588 357360 337660 357388
rect 319588 357348 319594 357360
rect 337654 357348 337660 357360
rect 337712 357348 337718 357400
rect 332410 354696 332416 354748
rect 332468 354736 332474 354748
rect 337654 354736 337660 354748
rect 332468 354708 337660 354736
rect 332468 354696 332474 354708
rect 337654 354696 337660 354708
rect 337712 354696 337718 354748
rect 330846 354084 330852 354136
rect 330904 354124 330910 354136
rect 337470 354124 337476 354136
rect 330904 354096 337476 354124
rect 330904 354084 330910 354096
rect 337470 354084 337476 354096
rect 337528 354084 337534 354136
rect 334618 353268 334624 353320
rect 334676 353308 334682 353320
rect 337746 353308 337752 353320
rect 334676 353280 337752 353308
rect 334676 353268 334682 353280
rect 337746 353268 337752 353280
rect 337804 353268 337810 353320
rect 329374 353200 329380 353252
rect 329432 353240 329438 353252
rect 337654 353240 337660 353252
rect 329432 353212 337660 353240
rect 329432 353200 329438 353212
rect 337654 353200 337660 353212
rect 337712 353200 337718 353252
rect 331858 351976 331864 352028
rect 331916 352016 331922 352028
rect 337286 352016 337292 352028
rect 331916 351988 337292 352016
rect 331916 351976 331922 351988
rect 337286 351976 337292 351988
rect 337344 351976 337350 352028
rect 323670 351908 323676 351960
rect 323728 351948 323734 351960
rect 336918 351948 336924 351960
rect 323728 351920 336924 351948
rect 323728 351908 323734 351920
rect 336918 351908 336924 351920
rect 336976 351908 336982 351960
rect 326522 351840 326528 351892
rect 326580 351880 326586 351892
rect 337654 351880 337660 351892
rect 326580 351852 337660 351880
rect 326580 351840 326586 351852
rect 337654 351840 337660 351852
rect 337712 351840 337718 351892
rect 330846 350548 330852 350600
rect 330904 350588 330910 350600
rect 337654 350588 337660 350600
rect 330904 350560 337660 350588
rect 330904 350548 330910 350560
rect 337654 350548 337660 350560
rect 337712 350548 337718 350600
rect 332318 350480 332324 350532
rect 332376 350520 332382 350532
rect 337746 350520 337752 350532
rect 332376 350492 337752 350520
rect 332376 350480 332382 350492
rect 337746 350480 337752 350492
rect 337804 350480 337810 350532
rect 328178 349120 328184 349172
rect 328236 349160 328242 349172
rect 337654 349160 337660 349172
rect 328236 349132 337660 349160
rect 328236 349120 328242 349132
rect 337654 349120 337660 349132
rect 337712 349120 337718 349172
rect 324038 349052 324044 349104
rect 324096 349092 324102 349104
rect 337746 349092 337752 349104
rect 324096 349064 337752 349092
rect 324096 349052 324102 349064
rect 337746 349052 337752 349064
rect 337804 349052 337810 349104
rect 334986 347284 334992 347336
rect 335044 347324 335050 347336
rect 337654 347324 337660 347336
rect 335044 347296 337660 347324
rect 335044 347284 335050 347296
rect 337654 347284 337660 347296
rect 337712 347284 337718 347336
rect 325418 347012 325424 347064
rect 325476 347052 325482 347064
rect 336918 347052 336924 347064
rect 325476 347024 336924 347052
rect 325476 347012 325482 347024
rect 336918 347012 336924 347024
rect 336976 347012 336982 347064
rect 325510 346400 325516 346452
rect 325568 346440 325574 346452
rect 337470 346440 337476 346452
rect 325568 346412 337476 346440
rect 325568 346400 325574 346412
rect 337470 346400 337476 346412
rect 337528 346400 337534 346452
rect 330754 346332 330760 346384
rect 330812 346372 330818 346384
rect 337654 346372 337660 346384
rect 330812 346344 337660 346372
rect 330812 346332 330818 346344
rect 337654 346332 337660 346344
rect 337712 346332 337718 346384
rect 334986 345040 334992 345092
rect 335044 345080 335050 345092
rect 337654 345080 337660 345092
rect 335044 345052 337660 345080
rect 335044 345040 335050 345052
rect 337654 345040 337660 345052
rect 337712 345040 337718 345092
rect 318058 344972 318064 345024
rect 318116 345012 318122 345024
rect 337746 345012 337752 345024
rect 318116 344984 337752 345012
rect 318116 344972 318122 344984
rect 337746 344972 337752 344984
rect 337804 344972 337810 345024
rect 324038 343612 324044 343664
rect 324096 343652 324102 343664
rect 337654 343652 337660 343664
rect 324096 343624 337660 343652
rect 324096 343612 324102 343624
rect 337654 343612 337660 343624
rect 337712 343612 337718 343664
rect 333330 343544 333336 343596
rect 333388 343584 333394 343596
rect 337562 343584 337568 343596
rect 333388 343556 337568 343584
rect 333388 343544 333394 343556
rect 337562 343544 337568 343556
rect 337620 343544 337626 343596
rect 329282 343476 329288 343528
rect 329340 343516 329346 343528
rect 337746 343516 337752 343528
rect 329340 343488 337752 343516
rect 329340 343476 329346 343488
rect 337746 343476 337752 343488
rect 337804 343476 337810 343528
rect 336274 342660 336280 342712
rect 336332 342700 336338 342712
rect 336734 342700 336740 342712
rect 336332 342672 336740 342700
rect 336332 342660 336338 342672
rect 336734 342660 336740 342672
rect 336792 342660 336798 342712
rect 322658 342252 322664 342304
rect 322716 342292 322722 342304
rect 337654 342292 337660 342304
rect 322716 342264 337660 342292
rect 322716 342252 322722 342264
rect 337654 342252 337660 342264
rect 337712 342252 337718 342304
rect 333330 339464 333336 339516
rect 333388 339504 333394 339516
rect 337286 339504 337292 339516
rect 333388 339476 337292 339504
rect 333388 339464 333394 339476
rect 337286 339464 337292 339476
rect 337344 339464 337350 339516
rect 332226 339396 332232 339448
rect 332284 339436 332290 339448
rect 337562 339436 337568 339448
rect 332284 339408 337568 339436
rect 332284 339396 332290 339408
rect 337562 339396 337568 339408
rect 337620 339396 337626 339448
rect 332318 338104 332324 338156
rect 332376 338144 332382 338156
rect 337286 338144 337292 338156
rect 332376 338116 337292 338144
rect 332376 338104 332382 338116
rect 337286 338104 337292 338116
rect 337344 338104 337350 338156
rect 326430 338036 326436 338088
rect 326488 338076 326494 338088
rect 337654 338076 337660 338088
rect 326488 338048 337660 338076
rect 326488 338036 326494 338048
rect 337654 338036 337660 338048
rect 337712 338036 337718 338088
rect 326522 336744 326528 336796
rect 326580 336784 326586 336796
rect 337746 336784 337752 336796
rect 326580 336756 337752 336784
rect 326580 336744 326586 336756
rect 337746 336744 337752 336756
rect 337804 336744 337810 336796
rect 321278 336676 321284 336728
rect 321336 336716 321342 336728
rect 337654 336716 337660 336728
rect 321336 336688 337660 336716
rect 321336 336676 321342 336688
rect 337654 336676 337660 336688
rect 337712 336676 337718 336728
rect 330754 335316 330760 335368
rect 330812 335356 330818 335368
rect 337838 335356 337844 335368
rect 330812 335328 337844 335356
rect 330812 335316 330818 335328
rect 337838 335316 337844 335328
rect 337896 335316 337902 335368
rect 323946 335248 323952 335300
rect 324004 335288 324010 335300
rect 337746 335288 337752 335300
rect 324004 335260 337752 335288
rect 324004 335248 324010 335260
rect 337746 335248 337752 335260
rect 337804 335248 337810 335300
rect 321278 333956 321284 334008
rect 321336 333996 321342 334008
rect 337562 333996 337568 334008
rect 321336 333968 337568 333996
rect 321336 333956 321342 333968
rect 337562 333956 337568 333968
rect 337620 333956 337626 334008
rect 323854 333208 323860 333260
rect 323912 333248 323918 333260
rect 337838 333248 337844 333260
rect 323912 333220 337844 333248
rect 323912 333208 323918 333220
rect 337838 333208 337844 333220
rect 337896 333208 337902 333260
rect 329374 332664 329380 332716
rect 329432 332704 329438 332716
rect 337654 332704 337660 332716
rect 329432 332676 337660 332704
rect 329432 332664 329438 332676
rect 337654 332664 337660 332676
rect 337712 332664 337718 332716
rect 323946 332596 323952 332648
rect 324004 332636 324010 332648
rect 337746 332636 337752 332648
rect 324004 332608 337752 332636
rect 324004 332596 324010 332608
rect 337746 332596 337752 332608
rect 337804 332596 337810 332648
rect 332134 332528 332140 332580
rect 332192 332568 332198 332580
rect 337654 332568 337660 332580
rect 332192 332540 337660 332568
rect 332192 332528 332198 332540
rect 337654 332528 337660 332540
rect 337712 332528 337718 332580
rect 160738 331168 160744 331220
rect 160796 331208 160802 331220
rect 161474 331208 161480 331220
rect 160796 331180 161480 331208
rect 160796 331168 160802 331180
rect 161474 331168 161480 331180
rect 161532 331208 161538 331220
rect 176654 331208 176660 331220
rect 161532 331180 176660 331208
rect 161532 331168 161538 331180
rect 176654 331168 176660 331180
rect 176712 331168 176718 331220
rect 322382 331168 322388 331220
rect 322440 331208 322446 331220
rect 337654 331208 337660 331220
rect 322440 331180 337660 331208
rect 322440 331168 322446 331180
rect 337654 331168 337660 331180
rect 337712 331168 337718 331220
rect 334894 331100 334900 331152
rect 334952 331140 334958 331152
rect 337562 331140 337568 331152
rect 334952 331112 337568 331140
rect 334952 331100 334958 331112
rect 337562 331100 337568 331112
rect 337620 331100 337626 331152
rect 335078 329808 335084 329860
rect 335136 329848 335142 329860
rect 337746 329848 337752 329860
rect 335136 329820 337752 329848
rect 335136 329808 335142 329820
rect 337746 329808 337752 329820
rect 337804 329808 337810 329860
rect 325234 329740 325240 329792
rect 325292 329780 325298 329792
rect 337654 329780 337660 329792
rect 325292 329752 337660 329780
rect 325292 329740 325298 329752
rect 337654 329740 337660 329752
rect 337712 329740 337718 329792
rect 332134 328448 332140 328500
rect 332192 328488 332198 328500
rect 337654 328488 337660 328500
rect 332192 328460 337660 328488
rect 332192 328448 332198 328460
rect 337654 328448 337660 328460
rect 337712 328448 337718 328500
rect 322382 327088 322388 327140
rect 322440 327128 322446 327140
rect 337102 327128 337108 327140
rect 322440 327100 337108 327128
rect 322440 327088 322446 327100
rect 337102 327088 337108 327100
rect 337160 327088 337166 327140
rect 330662 327020 330668 327072
rect 330720 327060 330726 327072
rect 337654 327060 337660 327072
rect 330720 327032 337660 327060
rect 330720 327020 330726 327032
rect 337654 327020 337660 327032
rect 337712 327020 337718 327072
rect 331122 325660 331128 325712
rect 331180 325700 331186 325712
rect 337654 325700 337660 325712
rect 331180 325672 337660 325700
rect 331180 325660 331186 325672
rect 337654 325660 337660 325672
rect 337712 325660 337718 325712
rect 321094 325592 321100 325644
rect 321152 325632 321158 325644
rect 337746 325632 337752 325644
rect 321152 325604 337752 325632
rect 321152 325592 321158 325604
rect 337746 325592 337752 325604
rect 337804 325592 337810 325644
rect 482278 325592 482284 325644
rect 482336 325632 482342 325644
rect 580166 325632 580172 325644
rect 482336 325604 580172 325632
rect 482336 325592 482342 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 318518 324300 318524 324352
rect 318576 324340 318582 324352
rect 337654 324340 337660 324352
rect 318576 324312 337660 324340
rect 318576 324300 318582 324312
rect 337654 324300 337660 324312
rect 337712 324300 337718 324352
rect 329282 322940 329288 322992
rect 329340 322980 329346 322992
rect 337654 322980 337660 322992
rect 329340 322952 337660 322980
rect 329340 322940 329346 322952
rect 337654 322940 337660 322952
rect 337712 322940 337718 322992
rect 156782 322396 156788 322448
rect 156840 322436 156846 322448
rect 337654 322436 337660 322448
rect 156840 322408 337660 322436
rect 156840 322396 156846 322408
rect 337654 322396 337660 322408
rect 337712 322396 337718 322448
rect 278682 322192 278688 322244
rect 278740 322232 278746 322244
rect 336458 322232 336464 322244
rect 278740 322204 336464 322232
rect 278740 322192 278746 322204
rect 336458 322192 336464 322204
rect 336516 322192 336522 322244
rect 179506 321784 179512 321836
rect 179564 321824 179570 321836
rect 223482 321824 223488 321836
rect 179564 321796 223488 321824
rect 179564 321784 179570 321796
rect 223482 321784 223488 321796
rect 223540 321784 223546 321836
rect 179414 321716 179420 321768
rect 179472 321756 179478 321768
rect 226334 321756 226340 321768
rect 179472 321728 226340 321756
rect 179472 321716 179478 321728
rect 226334 321716 226340 321728
rect 226392 321716 226398 321768
rect 179693 321691 179751 321697
rect 179693 321688 179705 321691
rect 178052 321660 179705 321688
rect 51074 321580 51080 321632
rect 51132 321620 51138 321632
rect 177945 321623 178003 321629
rect 177945 321620 177957 321623
rect 51132 321592 177957 321620
rect 51132 321580 51138 321592
rect 177945 321589 177957 321592
rect 177991 321589 178003 321623
rect 177945 321583 178003 321589
rect 62114 321512 62120 321564
rect 62172 321552 62178 321564
rect 62758 321552 62764 321564
rect 62172 321524 62764 321552
rect 62172 321512 62178 321524
rect 62758 321512 62764 321524
rect 62816 321552 62822 321564
rect 178052 321552 178080 321660
rect 179693 321657 179705 321660
rect 179739 321657 179751 321691
rect 179693 321651 179751 321657
rect 179782 321648 179788 321700
rect 179840 321688 179846 321700
rect 228634 321688 228640 321700
rect 179840 321660 228640 321688
rect 179840 321648 179846 321660
rect 228634 321648 228640 321660
rect 228692 321688 228698 321700
rect 229002 321688 229008 321700
rect 228692 321660 229008 321688
rect 228692 321648 228698 321660
rect 229002 321648 229008 321660
rect 229060 321648 229066 321700
rect 178129 321623 178187 321629
rect 178129 321589 178141 321623
rect 178175 321620 178187 321623
rect 204346 321620 204352 321632
rect 178175 321592 204352 321620
rect 178175 321589 178187 321592
rect 178129 321583 178187 321589
rect 204346 321580 204352 321592
rect 204404 321580 204410 321632
rect 231762 321580 231768 321632
rect 231820 321620 231826 321632
rect 337746 321620 337752 321632
rect 231820 321592 337752 321620
rect 231820 321580 231826 321592
rect 337746 321580 337752 321592
rect 337804 321580 337810 321632
rect 62816 321524 178080 321552
rect 179693 321555 179751 321561
rect 62816 321512 62822 321524
rect 179693 321521 179705 321555
rect 179739 321552 179751 321555
rect 180058 321552 180064 321564
rect 179739 321524 180064 321552
rect 179739 321521 179751 321524
rect 179693 321515 179751 321521
rect 180058 321512 180064 321524
rect 180116 321552 180122 321564
rect 185765 321555 185823 321561
rect 185765 321552 185777 321555
rect 180116 321524 185777 321552
rect 180116 321512 180122 321524
rect 185765 321521 185777 321524
rect 185811 321521 185823 321555
rect 185765 321515 185823 321521
rect 327902 321512 327908 321564
rect 327960 321552 327966 321564
rect 336918 321552 336924 321564
rect 327960 321524 336924 321552
rect 327960 321512 327966 321524
rect 336918 321512 336924 321524
rect 336976 321512 336982 321564
rect 71682 321444 71688 321496
rect 71740 321484 71746 321496
rect 337654 321484 337660 321496
rect 71740 321456 337660 321484
rect 71740 321444 71746 321456
rect 337654 321444 337660 321456
rect 337712 321444 337718 321496
rect 63494 321376 63500 321428
rect 63552 321416 63558 321428
rect 63862 321416 63868 321428
rect 63552 321388 63868 321416
rect 63552 321376 63558 321388
rect 63862 321376 63868 321388
rect 63920 321416 63926 321428
rect 177209 321419 177267 321425
rect 177209 321416 177221 321419
rect 63920 321388 177221 321416
rect 63920 321376 63926 321388
rect 177209 321385 177221 321388
rect 177255 321385 177267 321419
rect 177209 321379 177267 321385
rect 178218 321376 178224 321428
rect 178276 321416 178282 321428
rect 179322 321416 179328 321428
rect 178276 321388 179328 321416
rect 178276 321376 178282 321388
rect 179322 321376 179328 321388
rect 179380 321416 179386 321428
rect 219434 321416 219440 321428
rect 179380 321388 219440 321416
rect 179380 321376 179386 321388
rect 219434 321376 219440 321388
rect 219492 321416 219498 321428
rect 220630 321416 220636 321428
rect 219492 321388 220636 321416
rect 219492 321376 219498 321388
rect 220630 321376 220636 321388
rect 220688 321376 220694 321428
rect 246942 321376 246948 321428
rect 247000 321416 247006 321428
rect 326522 321416 326528 321428
rect 247000 321388 326528 321416
rect 247000 321376 247006 321388
rect 326522 321376 326528 321388
rect 326580 321376 326586 321428
rect 177025 321351 177083 321357
rect 177025 321317 177037 321351
rect 177071 321348 177083 321351
rect 179138 321348 179144 321360
rect 177071 321320 179144 321348
rect 177071 321317 177083 321320
rect 177025 321311 177083 321317
rect 179138 321308 179144 321320
rect 179196 321348 179202 321360
rect 220446 321348 220452 321360
rect 179196 321320 220452 321348
rect 179196 321308 179202 321320
rect 220446 321308 220452 321320
rect 220504 321308 220510 321360
rect 253842 321308 253848 321360
rect 253900 321348 253906 321360
rect 334986 321348 334992 321360
rect 253900 321320 334992 321348
rect 253900 321308 253906 321320
rect 334986 321308 334992 321320
rect 335044 321308 335050 321360
rect 178586 321240 178592 321292
rect 178644 321280 178650 321292
rect 203150 321280 203156 321292
rect 178644 321252 203156 321280
rect 178644 321240 178650 321252
rect 203150 321240 203156 321252
rect 203208 321240 203214 321292
rect 241422 321240 241428 321292
rect 241480 321280 241486 321292
rect 323946 321280 323952 321292
rect 241480 321252 323952 321280
rect 241480 321240 241486 321252
rect 323946 321240 323952 321252
rect 324004 321240 324010 321292
rect 117222 321172 117228 321224
rect 117280 321212 117286 321224
rect 329466 321212 329472 321224
rect 117280 321184 329472 321212
rect 117280 321172 117286 321184
rect 329466 321172 329472 321184
rect 329524 321172 329530 321224
rect 89622 321104 89628 321156
rect 89680 321144 89686 321156
rect 332318 321144 332324 321156
rect 89680 321116 332324 321144
rect 89680 321104 89686 321116
rect 332318 321104 332324 321116
rect 332376 321104 332382 321156
rect 86862 321036 86868 321088
rect 86920 321076 86926 321088
rect 330754 321076 330760 321088
rect 86920 321048 330760 321076
rect 86920 321036 86926 321048
rect 330754 321036 330760 321048
rect 330812 321036 330818 321088
rect 84102 320968 84108 321020
rect 84160 321008 84166 321020
rect 329374 321008 329380 321020
rect 84160 320980 329380 321008
rect 84160 320968 84166 320980
rect 329374 320968 329380 320980
rect 329432 320968 329438 321020
rect 77202 320900 77208 320952
rect 77260 320940 77266 320952
rect 331122 320940 331128 320952
rect 77260 320912 331128 320940
rect 77260 320900 77266 320912
rect 331122 320900 331128 320912
rect 331180 320900 331186 320952
rect 81342 320832 81348 320884
rect 81400 320872 81406 320884
rect 336182 320872 336188 320884
rect 81400 320844 336188 320872
rect 81400 320832 81406 320844
rect 336182 320832 336188 320844
rect 336240 320832 336246 320884
rect 60826 320764 60832 320816
rect 60884 320804 60890 320816
rect 177025 320807 177083 320813
rect 177025 320804 177037 320807
rect 60884 320776 177037 320804
rect 60884 320764 60890 320776
rect 177025 320773 177037 320776
rect 177071 320773 177083 320807
rect 177025 320767 177083 320773
rect 178034 320764 178040 320816
rect 178092 320804 178098 320816
rect 179230 320804 179236 320816
rect 178092 320776 179236 320804
rect 178092 320764 178098 320776
rect 179230 320764 179236 320776
rect 179288 320804 179294 320816
rect 211062 320804 211068 320816
rect 179288 320776 211068 320804
rect 179288 320764 179294 320776
rect 211062 320764 211068 320776
rect 211120 320764 211126 320816
rect 143350 320696 143356 320748
rect 143408 320736 143414 320748
rect 232038 320736 232044 320748
rect 143408 320708 232044 320736
rect 143408 320696 143414 320708
rect 232038 320696 232044 320708
rect 232096 320696 232102 320748
rect 143258 320628 143264 320680
rect 143316 320668 143322 320680
rect 233878 320668 233884 320680
rect 143316 320640 233884 320668
rect 143316 320628 143322 320640
rect 233878 320628 233884 320640
rect 233936 320628 233942 320680
rect 66162 320560 66168 320612
rect 66220 320600 66226 320612
rect 179414 320600 179420 320612
rect 66220 320572 179420 320600
rect 66220 320560 66226 320572
rect 179414 320560 179420 320572
rect 179472 320560 179478 320612
rect 179506 320560 179512 320612
rect 179564 320600 179570 320612
rect 215110 320600 215116 320612
rect 179564 320572 215116 320600
rect 179564 320560 179570 320572
rect 215110 320560 215116 320572
rect 215168 320560 215174 320612
rect 19978 320492 19984 320544
rect 20036 320532 20042 320544
rect 63494 320532 63500 320544
rect 20036 320504 63500 320532
rect 20036 320492 20042 320504
rect 63494 320492 63500 320504
rect 63552 320492 63558 320544
rect 176933 320535 176991 320541
rect 176933 320501 176945 320535
rect 176979 320532 176991 320535
rect 179046 320532 179052 320544
rect 176979 320504 179052 320532
rect 176979 320501 176991 320504
rect 176933 320495 176991 320501
rect 179046 320492 179052 320504
rect 179104 320532 179110 320544
rect 216398 320532 216404 320544
rect 179104 320504 216404 320532
rect 179104 320492 179110 320504
rect 216398 320492 216404 320504
rect 216456 320492 216462 320544
rect 19242 320424 19248 320476
rect 19300 320464 19306 320476
rect 62114 320464 62120 320476
rect 19300 320436 62120 320464
rect 19300 320424 19306 320436
rect 62114 320424 62120 320436
rect 62172 320424 62178 320476
rect 178126 320424 178132 320476
rect 178184 320464 178190 320476
rect 178770 320464 178776 320476
rect 178184 320436 178776 320464
rect 178184 320424 178190 320436
rect 178770 320424 178776 320436
rect 178828 320464 178834 320476
rect 216674 320464 216680 320476
rect 178828 320436 216680 320464
rect 178828 320424 178834 320436
rect 216674 320424 216680 320436
rect 216732 320424 216738 320476
rect 177209 320399 177267 320405
rect 177209 320365 177221 320399
rect 177255 320396 177267 320399
rect 179966 320396 179972 320408
rect 177255 320368 179972 320396
rect 177255 320365 177267 320368
rect 177209 320359 177267 320365
rect 179966 320356 179972 320368
rect 180024 320396 180030 320408
rect 185581 320399 185639 320405
rect 185581 320396 185593 320399
rect 180024 320368 185593 320396
rect 180024 320356 180030 320368
rect 185581 320365 185593 320368
rect 185627 320365 185639 320399
rect 185581 320359 185639 320365
rect 185673 320399 185731 320405
rect 185673 320365 185685 320399
rect 185719 320396 185731 320399
rect 218054 320396 218060 320408
rect 185719 320368 218060 320396
rect 185719 320365 185731 320368
rect 185673 320359 185731 320365
rect 218054 320356 218060 320368
rect 218112 320356 218118 320408
rect 60734 320288 60740 320340
rect 60792 320328 60798 320340
rect 178218 320328 178224 320340
rect 60792 320300 178224 320328
rect 60792 320288 60798 320300
rect 178218 320288 178224 320300
rect 178276 320288 178282 320340
rect 179414 320288 179420 320340
rect 179472 320328 179478 320340
rect 179874 320328 179880 320340
rect 179472 320300 179880 320328
rect 179472 320288 179478 320300
rect 179874 320288 179880 320300
rect 179932 320328 179938 320340
rect 202782 320328 202788 320340
rect 179932 320300 202788 320328
rect 179932 320288 179938 320300
rect 202782 320288 202788 320300
rect 202840 320288 202846 320340
rect 56594 320220 56600 320272
rect 56652 320260 56658 320272
rect 176933 320263 176991 320269
rect 176933 320260 176945 320263
rect 56652 320232 176945 320260
rect 56652 320220 56658 320232
rect 176933 320229 176945 320232
rect 176979 320229 176991 320263
rect 176933 320223 176991 320229
rect 177945 320263 178003 320269
rect 177945 320229 177957 320263
rect 177991 320260 178003 320263
rect 181073 320263 181131 320269
rect 181073 320260 181085 320263
rect 177991 320232 181085 320260
rect 177991 320229 178003 320232
rect 177945 320223 178003 320229
rect 181073 320229 181085 320232
rect 181119 320229 181131 320263
rect 185489 320263 185547 320269
rect 185489 320260 185501 320263
rect 181073 320223 181131 320229
rect 181180 320232 185501 320260
rect 19150 320152 19156 320204
rect 19208 320192 19214 320204
rect 65334 320192 65340 320204
rect 19208 320164 65340 320192
rect 19208 320152 19214 320164
rect 65334 320152 65340 320164
rect 65392 320192 65398 320204
rect 66162 320192 66168 320204
rect 65392 320164 66168 320192
rect 65392 320152 65398 320164
rect 66162 320152 66168 320164
rect 66220 320152 66226 320204
rect 176856 320164 180104 320192
rect 18874 320084 18880 320136
rect 18932 320124 18938 320136
rect 44174 320124 44180 320136
rect 18932 320096 44180 320124
rect 18932 320084 18938 320096
rect 44174 320084 44180 320096
rect 44232 320124 44238 320136
rect 51074 320124 51080 320136
rect 44232 320096 51080 320124
rect 44232 320084 44238 320096
rect 51074 320084 51080 320096
rect 51132 320084 51138 320136
rect 79226 320084 79232 320136
rect 79284 320124 79290 320136
rect 157334 320124 157340 320136
rect 79284 320096 157340 320124
rect 79284 320084 79290 320096
rect 157334 320084 157340 320096
rect 157392 320084 157398 320136
rect 19058 320016 19064 320068
rect 19116 320056 19122 320068
rect 50154 320056 50160 320068
rect 19116 320028 50160 320056
rect 19116 320016 19122 320028
rect 50154 320016 50160 320028
rect 50212 320016 50218 320068
rect 50249 320059 50307 320065
rect 50249 320025 50261 320059
rect 50295 320056 50307 320059
rect 51258 320056 51264 320068
rect 50295 320028 51264 320056
rect 50295 320025 50307 320028
rect 50249 320019 50307 320025
rect 51258 320016 51264 320028
rect 51316 320056 51322 320068
rect 60001 320059 60059 320065
rect 60001 320056 60013 320059
rect 51316 320028 60013 320056
rect 51316 320016 51322 320028
rect 60001 320025 60013 320028
rect 60047 320025 60059 320059
rect 60001 320019 60059 320025
rect 77294 320016 77300 320068
rect 77352 320056 77358 320068
rect 176378 320056 176384 320068
rect 77352 320028 176384 320056
rect 77352 320016 77358 320028
rect 176378 320016 176384 320028
rect 176436 320056 176442 320068
rect 176856 320056 176884 320164
rect 177942 320124 177948 320136
rect 176436 320028 176884 320056
rect 176948 320096 177948 320124
rect 176436 320016 176442 320028
rect 18414 319948 18420 320000
rect 18472 319988 18478 320000
rect 59354 319988 59360 320000
rect 18472 319960 59360 319988
rect 18472 319948 18478 319960
rect 59354 319948 59360 319960
rect 59412 319948 59418 320000
rect 78674 319948 78680 320000
rect 78732 319988 78738 320000
rect 176948 319988 176976 320096
rect 177942 320084 177948 320096
rect 178000 320124 178006 320136
rect 179969 320127 180027 320133
rect 179969 320124 179981 320127
rect 178000 320096 179981 320124
rect 178000 320084 178006 320096
rect 179969 320093 179981 320096
rect 180015 320093 180027 320127
rect 180076 320124 180104 320164
rect 180150 320152 180156 320204
rect 180208 320192 180214 320204
rect 181180 320192 181208 320232
rect 185489 320229 185501 320232
rect 185535 320229 185547 320263
rect 185489 320223 185547 320229
rect 185581 320263 185639 320269
rect 185581 320229 185593 320263
rect 185627 320260 185639 320263
rect 204898 320260 204904 320272
rect 185627 320232 204904 320260
rect 185627 320229 185639 320232
rect 185581 320223 185639 320229
rect 204898 320220 204904 320232
rect 204956 320220 204962 320272
rect 180208 320164 181208 320192
rect 181257 320195 181315 320201
rect 180208 320152 180214 320164
rect 181257 320161 181269 320195
rect 181303 320192 181315 320195
rect 185765 320195 185823 320201
rect 181303 320164 185716 320192
rect 181303 320161 181315 320164
rect 181257 320155 181315 320161
rect 185688 320124 185716 320164
rect 185765 320161 185777 320195
rect 185811 320192 185823 320195
rect 208394 320192 208400 320204
rect 185811 320164 208400 320192
rect 185811 320161 185823 320164
rect 185765 320155 185823 320161
rect 208394 320152 208400 320164
rect 208452 320152 208458 320204
rect 200758 320124 200764 320136
rect 180076 320096 185624 320124
rect 185688 320096 200764 320124
rect 179969 320087 180027 320093
rect 179782 320056 179788 320068
rect 78732 319960 176976 319988
rect 177040 320028 179788 320056
rect 78732 319948 78738 319960
rect 19518 319880 19524 319932
rect 19576 319920 19582 319932
rect 75730 319920 75736 319932
rect 19576 319892 75736 319920
rect 19576 319880 19582 319892
rect 75730 319880 75736 319892
rect 75788 319920 75794 319932
rect 177040 319920 177068 320028
rect 179782 320016 179788 320028
rect 179840 320016 179846 320068
rect 179877 320059 179935 320065
rect 179877 320025 179889 320059
rect 179923 320056 179935 320059
rect 185489 320059 185547 320065
rect 185489 320056 185501 320059
rect 179923 320028 185501 320056
rect 179923 320025 179935 320028
rect 179877 320019 179935 320025
rect 185489 320025 185501 320028
rect 185535 320025 185547 320059
rect 185596 320056 185624 320096
rect 200758 320084 200764 320096
rect 200816 320084 200822 320136
rect 204898 320084 204904 320136
rect 204956 320124 204962 320136
rect 224126 320124 224132 320136
rect 204956 320096 224132 320124
rect 204956 320084 204962 320096
rect 224126 320084 224132 320096
rect 224184 320084 224190 320136
rect 334802 320084 334808 320136
rect 334860 320124 334866 320136
rect 337654 320124 337660 320136
rect 334860 320096 337660 320124
rect 334860 320084 334866 320096
rect 337654 320084 337660 320096
rect 337712 320084 337718 320136
rect 236638 320056 236644 320068
rect 185596 320028 236644 320056
rect 185489 320019 185547 320025
rect 236638 320016 236644 320028
rect 236696 320016 236702 320068
rect 178126 319948 178132 320000
rect 178184 319988 178190 320000
rect 180061 319991 180119 319997
rect 178184 319960 179828 319988
rect 178184 319948 178190 319960
rect 179690 319920 179696 319932
rect 75788 319892 177068 319920
rect 177960 319892 179696 319920
rect 75788 319880 75794 319892
rect 19886 319812 19892 319864
rect 19944 319852 19950 319864
rect 66438 319852 66444 319864
rect 19944 319824 66444 319852
rect 19944 319812 19950 319824
rect 66438 319812 66444 319824
rect 66496 319812 66502 319864
rect 74626 319812 74632 319864
rect 74684 319852 74690 319864
rect 177960 319852 177988 319892
rect 179690 319880 179696 319892
rect 179748 319880 179754 319932
rect 74684 319824 177988 319852
rect 74684 319812 74690 319824
rect 178034 319812 178040 319864
rect 178092 319852 178098 319864
rect 179800 319852 179828 319960
rect 180061 319957 180073 319991
rect 180107 319988 180119 319991
rect 211798 319988 211804 320000
rect 180107 319960 211804 319988
rect 180107 319957 180119 319960
rect 180061 319951 180119 319957
rect 211798 319948 211804 319960
rect 211856 319948 211862 320000
rect 179877 319923 179935 319929
rect 179877 319889 179889 319923
rect 179923 319920 179935 319923
rect 185397 319923 185455 319929
rect 185397 319920 185409 319923
rect 179923 319892 185409 319920
rect 179923 319889 179935 319892
rect 179877 319883 179935 319889
rect 185397 319889 185409 319892
rect 185443 319889 185455 319923
rect 185397 319883 185455 319889
rect 185489 319923 185547 319929
rect 185489 319889 185501 319923
rect 185535 319920 185547 319923
rect 229554 319920 229560 319932
rect 185535 319892 229560 319920
rect 185535 319889 185547 319892
rect 185489 319883 185547 319889
rect 229554 319880 229560 319892
rect 229612 319880 229618 319932
rect 271782 319880 271788 319932
rect 271840 319920 271846 319932
rect 322566 319920 322572 319932
rect 271840 319892 322572 319920
rect 271840 319880 271846 319892
rect 322566 319880 322572 319892
rect 322624 319880 322630 319932
rect 178092 319824 179736 319852
rect 179800 319824 209774 319852
rect 178092 319812 178098 319824
rect 18138 319744 18144 319796
rect 18196 319784 18202 319796
rect 73338 319784 73344 319796
rect 18196 319756 73344 319784
rect 18196 319744 18202 319756
rect 73338 319744 73344 319756
rect 73396 319784 73402 319796
rect 179598 319784 179604 319796
rect 73396 319756 179604 319784
rect 73396 319744 73402 319756
rect 179598 319744 179604 319756
rect 179656 319744 179662 319796
rect 179708 319784 179736 319824
rect 185765 319787 185823 319793
rect 179708 319756 185716 319784
rect 19702 319676 19708 319728
rect 19760 319716 19766 319728
rect 68646 319716 68652 319728
rect 19760 319688 68652 319716
rect 19760 319676 19766 319688
rect 68646 319676 68652 319688
rect 68704 319676 68710 319728
rect 70394 319676 70400 319728
rect 70452 319716 70458 319728
rect 176470 319716 176476 319728
rect 70452 319688 176476 319716
rect 70452 319676 70458 319688
rect 176470 319676 176476 319688
rect 176528 319676 176534 319728
rect 176562 319676 176568 319728
rect 176620 319716 176626 319728
rect 177945 319719 178003 319725
rect 177945 319716 177957 319719
rect 176620 319688 177957 319716
rect 176620 319676 176626 319688
rect 177945 319685 177957 319688
rect 177991 319685 178003 319719
rect 178494 319716 178500 319728
rect 177945 319679 178003 319685
rect 178052 319688 178500 319716
rect 18230 319608 18236 319660
rect 18288 319648 18294 319660
rect 72142 319648 72148 319660
rect 18288 319620 72148 319648
rect 18288 319608 18294 319620
rect 72142 319608 72148 319620
rect 72200 319648 72206 319660
rect 178052 319648 178080 319688
rect 178494 319676 178500 319688
rect 178552 319716 178558 319728
rect 185688 319716 185716 319756
rect 185765 319753 185777 319787
rect 185811 319784 185823 319787
rect 204901 319787 204959 319793
rect 204901 319784 204913 319787
rect 185811 319756 204913 319784
rect 185811 319753 185823 319756
rect 185765 319747 185823 319753
rect 204901 319753 204913 319756
rect 204947 319753 204959 319787
rect 209746 319784 209774 319824
rect 211062 319812 211068 319864
rect 211120 319852 211126 319864
rect 221826 319852 221832 319864
rect 211120 319824 221832 319852
rect 211120 319812 211126 319824
rect 221826 319812 221832 319824
rect 221884 319852 221890 319864
rect 222102 319852 222108 319864
rect 221884 319824 222108 319852
rect 221884 319812 221890 319824
rect 222102 319812 222108 319824
rect 222160 319812 222166 319864
rect 277302 319812 277308 319864
rect 277360 319852 277366 319864
rect 333422 319852 333428 319864
rect 277360 319824 333428 319852
rect 277360 319812 277366 319824
rect 333422 319812 333428 319824
rect 333480 319812 333486 319864
rect 210418 319784 210424 319796
rect 209746 319756 210424 319784
rect 204901 319747 204959 319753
rect 210418 319744 210424 319756
rect 210476 319744 210482 319796
rect 269022 319744 269028 319796
rect 269080 319784 269086 319796
rect 329558 319784 329564 319796
rect 269080 319756 329564 319784
rect 269080 319744 269086 319756
rect 329558 319744 329564 319756
rect 329616 319744 329622 319796
rect 207290 319716 207296 319728
rect 178552 319688 185624 319716
rect 185688 319688 207296 319716
rect 178552 319676 178558 319688
rect 72200 319620 178080 319648
rect 72200 319608 72206 319620
rect 179414 319608 179420 319660
rect 179472 319648 179478 319660
rect 180518 319648 180524 319660
rect 179472 319620 180524 319648
rect 179472 319608 179478 319620
rect 180518 319608 180524 319620
rect 180576 319648 180582 319660
rect 185596 319648 185624 319688
rect 207290 319676 207296 319688
rect 207348 319676 207354 319728
rect 208394 319676 208400 319728
rect 208452 319716 208458 319728
rect 222838 319716 222844 319728
rect 208452 319688 222844 319716
rect 208452 319676 208458 319688
rect 222838 319676 222844 319688
rect 222896 319676 222902 319728
rect 274542 319676 274548 319728
rect 274600 319716 274606 319728
rect 335170 319716 335176 319728
rect 274600 319688 335176 319716
rect 274600 319676 274606 319688
rect 335170 319676 335176 319688
rect 335228 319676 335234 319728
rect 231854 319648 231860 319660
rect 180576 319620 185072 319648
rect 185596 319620 231860 319648
rect 180576 319608 180582 319620
rect 17310 319540 17316 319592
rect 17368 319580 17374 319592
rect 71130 319580 71136 319592
rect 17368 319552 71136 319580
rect 17368 319540 17374 319552
rect 71130 319540 71136 319552
rect 71188 319580 71194 319592
rect 179506 319580 179512 319592
rect 71188 319552 179512 319580
rect 71188 319540 71194 319552
rect 179506 319540 179512 319552
rect 179564 319580 179570 319592
rect 185044 319580 185072 319620
rect 231854 319608 231860 319620
rect 231912 319608 231918 319660
rect 264882 319608 264888 319660
rect 264940 319648 264946 319660
rect 332410 319648 332416 319660
rect 264940 319620 332416 319648
rect 264940 319608 264946 319620
rect 332410 319608 332416 319620
rect 332468 319608 332474 319660
rect 213178 319580 213184 319592
rect 179564 319552 184980 319580
rect 185044 319552 213184 319580
rect 179564 319540 179570 319552
rect 18598 319472 18604 319524
rect 18656 319512 18662 319524
rect 52362 319512 52368 319524
rect 18656 319484 52368 319512
rect 18656 319472 18662 319484
rect 52362 319472 52368 319484
rect 52420 319512 52426 319524
rect 178586 319512 178592 319524
rect 52420 319484 178592 319512
rect 52420 319472 52426 319484
rect 178586 319472 178592 319484
rect 178644 319512 178650 319524
rect 179877 319515 179935 319521
rect 179877 319512 179889 319515
rect 178644 319484 179889 319512
rect 178644 319472 178650 319484
rect 179877 319481 179889 319484
rect 179923 319481 179935 319515
rect 179877 319475 179935 319481
rect 179969 319515 180027 319521
rect 179969 319481 179981 319515
rect 180015 319512 180027 319515
rect 181993 319515 182051 319521
rect 181993 319512 182005 319515
rect 180015 319484 182005 319512
rect 180015 319481 180027 319484
rect 179969 319475 180027 319481
rect 181993 319481 182005 319484
rect 182039 319481 182051 319515
rect 184952 319512 184980 319552
rect 213178 319540 213184 319552
rect 213236 319540 213242 319592
rect 233878 319540 233884 319592
rect 233936 319580 233942 319592
rect 303062 319580 303068 319592
rect 233936 319552 303068 319580
rect 233936 319540 233942 319552
rect 303062 319540 303068 319552
rect 303120 319540 303126 319592
rect 231210 319512 231216 319524
rect 184952 319484 231216 319512
rect 181993 319475 182051 319481
rect 231210 319472 231216 319484
rect 231268 319512 231274 319524
rect 231670 319512 231676 319524
rect 231268 319484 231676 319512
rect 231268 319472 231274 319484
rect 231670 319472 231676 319484
rect 231728 319472 231734 319524
rect 232038 319472 232044 319524
rect 232096 319512 232102 319524
rect 302878 319512 302884 319524
rect 232096 319484 302884 319512
rect 232096 319472 232102 319484
rect 302878 319472 302884 319484
rect 302936 319472 302942 319524
rect 19610 319404 19616 319456
rect 19668 319444 19674 319456
rect 53466 319444 53472 319456
rect 19668 319416 53472 319444
rect 19668 319404 19674 319416
rect 53466 319404 53472 319416
rect 53524 319444 53530 319456
rect 179414 319444 179420 319456
rect 53524 319416 179420 319444
rect 53524 319404 53530 319416
rect 179414 319404 179420 319416
rect 179472 319404 179478 319456
rect 179598 319404 179604 319456
rect 179656 319444 179662 319456
rect 233878 319444 233884 319456
rect 179656 319416 233884 319444
rect 179656 319404 179662 319416
rect 233878 319404 233884 319416
rect 233936 319404 233942 319456
rect 256602 319404 256608 319456
rect 256660 319444 256666 319456
rect 336366 319444 336372 319456
rect 256660 319416 336372 319444
rect 256660 319404 256666 319416
rect 336366 319404 336372 319416
rect 336424 319404 336430 319456
rect 18966 319336 18972 319388
rect 19024 319376 19030 319388
rect 59906 319376 59912 319388
rect 19024 319348 59912 319376
rect 19024 319336 19030 319348
rect 59906 319336 59912 319348
rect 59964 319336 59970 319388
rect 60001 319379 60059 319385
rect 60001 319345 60013 319379
rect 60047 319376 60059 319379
rect 178862 319376 178868 319388
rect 60047 319348 178868 319376
rect 60047 319345 60059 319348
rect 60001 319339 60059 319345
rect 178862 319336 178868 319348
rect 178920 319376 178926 319388
rect 178920 319348 179644 319376
rect 178920 319336 178926 319348
rect 18506 319268 18512 319320
rect 18564 319308 18570 319320
rect 50065 319311 50123 319317
rect 50065 319308 50077 319311
rect 18564 319280 50077 319308
rect 18564 319268 18570 319280
rect 50065 319277 50077 319280
rect 50111 319277 50123 319311
rect 50065 319271 50123 319277
rect 50154 319268 50160 319320
rect 50212 319308 50218 319320
rect 178126 319308 178132 319320
rect 50212 319280 178132 319308
rect 50212 319268 50218 319280
rect 178126 319268 178132 319280
rect 178184 319308 178190 319320
rect 178770 319308 178776 319320
rect 178184 319280 178776 319308
rect 178184 319268 178190 319280
rect 178770 319268 178776 319280
rect 178828 319268 178834 319320
rect 179509 319311 179567 319317
rect 179509 319308 179521 319311
rect 179340 319280 179521 319308
rect 40678 319200 40684 319252
rect 40736 319240 40742 319252
rect 176286 319240 176292 319252
rect 40736 319212 176292 319240
rect 40736 319200 40742 319212
rect 176286 319200 176292 319212
rect 176344 319200 176350 319252
rect 176470 319200 176476 319252
rect 176528 319240 176534 319252
rect 179340 319240 179368 319280
rect 179509 319277 179521 319280
rect 179555 319277 179567 319311
rect 179616 319308 179644 319348
rect 179690 319336 179696 319388
rect 179748 319376 179754 319388
rect 234062 319376 234068 319388
rect 179748 319348 234068 319376
rect 179748 319336 179754 319348
rect 234062 319336 234068 319348
rect 234120 319336 234126 319388
rect 180061 319311 180119 319317
rect 180061 319308 180073 319311
rect 179616 319280 180073 319308
rect 179509 319271 179567 319277
rect 180061 319277 180073 319280
rect 180107 319277 180119 319311
rect 235258 319308 235264 319320
rect 180061 319271 180119 319277
rect 180766 319280 235264 319308
rect 176528 319212 179368 319240
rect 176528 319200 176534 319212
rect 179414 319200 179420 319252
rect 179472 319240 179478 319252
rect 179782 319240 179788 319252
rect 179472 319212 179788 319240
rect 179472 319200 179478 319212
rect 179782 319200 179788 319212
rect 179840 319240 179846 319252
rect 180766 319240 180794 319280
rect 235258 319268 235264 319280
rect 235316 319268 235322 319320
rect 179840 319212 180794 319240
rect 181993 319243 182051 319249
rect 179840 319200 179846 319212
rect 181993 319209 182005 319243
rect 182039 319240 182051 319243
rect 238018 319240 238024 319252
rect 182039 319212 238024 319240
rect 182039 319209 182051 319212
rect 181993 319203 182051 319209
rect 238018 319200 238024 319212
rect 238076 319200 238082 319252
rect 42058 319132 42064 319184
rect 42116 319172 42122 319184
rect 178678 319172 178684 319184
rect 42116 319144 178684 319172
rect 42116 319132 42122 319144
rect 178678 319132 178684 319144
rect 178736 319172 178742 319184
rect 201494 319172 201500 319184
rect 178736 319144 201500 319172
rect 178736 319132 178742 319144
rect 201494 319132 201500 319144
rect 201552 319172 201558 319184
rect 202138 319172 202144 319184
rect 201552 319144 202144 319172
rect 201552 319132 201558 319144
rect 202138 319132 202144 319144
rect 202196 319132 202202 319184
rect 202782 319132 202788 319184
rect 202840 319172 202846 319184
rect 225598 319172 225604 319184
rect 202840 319144 225604 319172
rect 202840 319132 202846 319144
rect 225598 319132 225604 319144
rect 225656 319132 225662 319184
rect 20070 319064 20076 319116
rect 20128 319104 20134 319116
rect 36078 319104 36084 319116
rect 20128 319076 36084 319104
rect 20128 319064 20134 319076
rect 36078 319064 36084 319076
rect 36136 319104 36142 319116
rect 196066 319104 196072 319116
rect 36136 319076 196072 319104
rect 36136 319064 36142 319076
rect 196066 319064 196072 319076
rect 196124 319064 196130 319116
rect 204901 319107 204959 319113
rect 204901 319073 204913 319107
rect 204947 319104 204959 319107
rect 211338 319104 211344 319116
rect 204947 319076 211344 319104
rect 204947 319073 204959 319076
rect 204901 319067 204959 319073
rect 211338 319064 211344 319076
rect 211396 319064 211402 319116
rect 37918 318996 37924 319048
rect 37976 319036 37982 319048
rect 197354 319036 197360 319048
rect 37976 319008 197360 319036
rect 37976 318996 37982 319008
rect 197354 318996 197360 319008
rect 197412 318996 197418 319048
rect 18782 318928 18788 318980
rect 18840 318968 18846 318980
rect 39574 318968 39580 318980
rect 18840 318940 39580 318968
rect 18840 318928 18846 318940
rect 39574 318928 39580 318940
rect 39632 318968 39638 318980
rect 198734 318968 198740 318980
rect 39632 318940 198740 318968
rect 39632 318928 39638 318940
rect 198734 318928 198740 318940
rect 198792 318928 198798 318980
rect 231670 318928 231676 318980
rect 231728 318968 231734 318980
rect 316770 318968 316776 318980
rect 231728 318940 316776 318968
rect 231728 318928 231734 318940
rect 316770 318928 316776 318940
rect 316828 318928 316834 318980
rect 36538 318860 36544 318912
rect 36596 318900 36602 318912
rect 195974 318900 195980 318912
rect 36596 318872 195980 318900
rect 36596 318860 36602 318872
rect 195974 318860 195980 318872
rect 196032 318860 196038 318912
rect 224126 318860 224132 318912
rect 224184 318900 224190 318912
rect 316678 318900 316684 318912
rect 224184 318872 316684 318900
rect 224184 318860 224190 318872
rect 316678 318860 316684 318872
rect 316736 318860 316742 318912
rect 18322 318792 18328 318844
rect 18380 318832 18386 318844
rect 45002 318832 45008 318844
rect 18380 318804 45008 318832
rect 18380 318792 18386 318804
rect 45002 318792 45008 318804
rect 45060 318832 45066 318844
rect 204254 318832 204260 318844
rect 45060 318804 204260 318832
rect 45060 318792 45066 318804
rect 204254 318792 204260 318804
rect 204312 318792 204318 318844
rect 228910 318792 228916 318844
rect 228968 318832 228974 318844
rect 337746 318832 337752 318844
rect 228968 318804 337752 318832
rect 228968 318792 228974 318804
rect 337746 318792 337752 318804
rect 337804 318792 337810 318844
rect 176286 318724 176292 318776
rect 176344 318764 176350 318776
rect 176562 318764 176568 318776
rect 176344 318736 176568 318764
rect 176344 318724 176350 318736
rect 176562 318724 176568 318736
rect 176620 318724 176626 318776
rect 281442 318724 281448 318776
rect 281500 318764 281506 318776
rect 326614 318764 326620 318776
rect 281500 318736 326620 318764
rect 281500 318724 281506 318736
rect 326614 318724 326620 318736
rect 326672 318724 326678 318776
rect 259362 318656 259368 318708
rect 259420 318696 259426 318708
rect 330846 318696 330852 318708
rect 259420 318668 330852 318696
rect 259420 318656 259426 318668
rect 330846 318656 330852 318668
rect 330904 318656 330910 318708
rect 251082 318588 251088 318640
rect 251140 318628 251146 318640
rect 322658 318628 322664 318640
rect 251140 318600 322664 318628
rect 251140 318588 251146 318600
rect 322658 318588 322664 318600
rect 322716 318588 322722 318640
rect 326338 318588 326344 318640
rect 326396 318628 326402 318640
rect 337654 318628 337660 318640
rect 326396 318600 337660 318628
rect 326396 318588 326402 318600
rect 337654 318588 337660 318600
rect 337712 318588 337718 318640
rect 249702 318520 249708 318572
rect 249760 318560 249766 318572
rect 333330 318560 333336 318572
rect 249760 318532 333336 318560
rect 249760 318520 249766 318532
rect 333330 318520 333336 318532
rect 333388 318520 333394 318572
rect 222102 318452 222108 318504
rect 222160 318492 222166 318504
rect 323854 318492 323860 318504
rect 222160 318464 323860 318492
rect 222160 318452 222166 318464
rect 323854 318452 323860 318464
rect 323912 318452 323918 318504
rect 207290 318384 207296 318436
rect 207348 318424 207354 318436
rect 330662 318424 330668 318436
rect 207348 318396 330668 318424
rect 207348 318384 207354 318396
rect 330662 318384 330668 318396
rect 330720 318384 330726 318436
rect 179598 318316 179604 318368
rect 179656 318356 179662 318368
rect 179782 318356 179788 318368
rect 179656 318328 179788 318356
rect 179656 318316 179662 318328
rect 179782 318316 179788 318328
rect 179840 318316 179846 318368
rect 203794 318316 203800 318368
rect 203852 318356 203858 318368
rect 334802 318356 334808 318368
rect 203852 318328 334808 318356
rect 203852 318316 203858 318328
rect 334802 318316 334808 318328
rect 334860 318316 334866 318368
rect 159358 318248 159364 318300
rect 159416 318288 159422 318300
rect 336182 318288 336188 318300
rect 159416 318260 336188 318288
rect 159416 318248 159422 318260
rect 336182 318248 336188 318260
rect 336240 318248 336246 318300
rect 99282 318180 99288 318232
rect 99340 318220 99346 318232
rect 328178 318220 328184 318232
rect 99340 318192 328184 318220
rect 99340 318180 99346 318192
rect 328178 318180 328184 318192
rect 328236 318180 328242 318232
rect 93762 318112 93768 318164
rect 93820 318152 93826 318164
rect 324038 318152 324044 318164
rect 93820 318124 324044 318152
rect 93820 318112 93826 318124
rect 324038 318112 324044 318124
rect 324096 318112 324102 318164
rect 91002 318044 91008 318096
rect 91060 318084 91066 318096
rect 336274 318084 336280 318096
rect 91060 318056 336280 318084
rect 91060 318044 91066 318056
rect 336274 318044 336280 318056
rect 336332 318044 336338 318096
rect 68922 317432 68928 317484
rect 68980 317472 68986 317484
rect 336918 317472 336924 317484
rect 68980 317444 336924 317472
rect 68980 317432 68986 317444
rect 336918 317432 336924 317444
rect 336976 317432 336982 317484
rect 156690 317364 156696 317416
rect 156748 317404 156754 317416
rect 337654 317404 337660 317416
rect 156748 317376 337660 317404
rect 156748 317364 156754 317376
rect 337654 317364 337660 317376
rect 337712 317364 337718 317416
rect 226242 316004 226248 316056
rect 226300 316044 226306 316056
rect 337562 316044 337568 316056
rect 226300 316016 337568 316044
rect 226300 316004 226306 316016
rect 337562 316004 337568 316016
rect 337620 316004 337626 316056
rect 329190 315936 329196 315988
rect 329248 315976 329254 315988
rect 337654 315976 337660 315988
rect 329248 315948 337660 315976
rect 329248 315936 329254 315948
rect 337654 315936 337660 315948
rect 337712 315936 337718 315988
rect 238662 315256 238668 315308
rect 238720 315296 238726 315308
rect 335078 315296 335084 315308
rect 238720 315268 335084 315296
rect 238720 315256 238726 315268
rect 335078 315256 335084 315268
rect 335136 315256 335142 315308
rect 223482 314712 223488 314764
rect 223540 314752 223546 314764
rect 337654 314752 337660 314764
rect 223540 314724 337660 314752
rect 223540 314712 223546 314724
rect 337654 314712 337660 314724
rect 337712 314712 337718 314764
rect 66162 314644 66168 314696
rect 66220 314684 66226 314696
rect 337746 314684 337752 314696
rect 66220 314656 337752 314684
rect 66220 314644 66226 314656
rect 337746 314644 337752 314656
rect 337804 314644 337810 314696
rect 156598 314576 156604 314628
rect 156656 314616 156662 314628
rect 337654 314616 337660 314628
rect 156656 314588 337660 314616
rect 156656 314576 156662 314588
rect 337654 314576 337660 314588
rect 337712 314576 337718 314628
rect 64782 313284 64788 313336
rect 64840 313324 64846 313336
rect 337654 313324 337660 313336
rect 64840 313296 337660 313324
rect 64840 313284 64846 313296
rect 337654 313284 337660 313296
rect 337712 313284 337718 313336
rect 325142 313216 325148 313268
rect 325200 313256 325206 313268
rect 337746 313256 337752 313268
rect 325200 313228 337752 313256
rect 325200 313216 325206 313228
rect 337746 313216 337752 313228
rect 337804 313216 337810 313268
rect 482370 313216 482376 313268
rect 482428 313256 482434 313268
rect 580166 313256 580172 313268
rect 482428 313228 580172 313256
rect 482428 313216 482434 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 219250 312536 219256 312588
rect 219308 312576 219314 312588
rect 327902 312576 327908 312588
rect 219308 312548 327908 312576
rect 219308 312536 219314 312548
rect 327902 312536 327908 312548
rect 327960 312536 327966 312588
rect 222102 311856 222108 311908
rect 222160 311896 222166 311908
rect 337746 311896 337752 311908
rect 222160 311868 337752 311896
rect 222160 311856 222166 311868
rect 337746 311856 337752 311868
rect 337804 311856 337810 311908
rect 178402 311788 178408 311840
rect 178460 311828 178466 311840
rect 337654 311828 337660 311840
rect 178460 311800 337660 311828
rect 178460 311788 178466 311800
rect 337654 311788 337660 311800
rect 337712 311788 337718 311840
rect 62022 310496 62028 310548
rect 62080 310536 62086 310548
rect 337654 310536 337660 310548
rect 62080 310508 337660 310536
rect 62080 310496 62086 310508
rect 337654 310496 337660 310508
rect 337712 310496 337718 310548
rect 332042 310428 332048 310480
rect 332100 310468 332106 310480
rect 337102 310468 337108 310480
rect 332100 310440 337108 310468
rect 332100 310428 332106 310440
rect 337102 310428 337108 310440
rect 337160 310428 337166 310480
rect 219342 309136 219348 309188
rect 219400 309176 219406 309188
rect 337654 309176 337660 309188
rect 219400 309148 337660 309176
rect 219400 309136 219406 309148
rect 337654 309136 337660 309148
rect 337712 309136 337718 309188
rect 173158 309068 173164 309120
rect 173216 309108 173222 309120
rect 337102 309108 337108 309120
rect 173216 309080 337108 309108
rect 173216 309068 173222 309080
rect 337102 309068 337108 309080
rect 337160 309068 337166 309120
rect 59262 307776 59268 307828
rect 59320 307816 59326 307828
rect 337654 307816 337660 307828
rect 59320 307788 337660 307816
rect 59320 307776 59326 307788
rect 337654 307776 337660 307788
rect 337712 307776 337718 307828
rect 170398 307708 170404 307760
rect 170456 307748 170462 307760
rect 337746 307748 337752 307760
rect 170456 307720 337752 307748
rect 170456 307708 170462 307720
rect 337746 307708 337752 307720
rect 337804 307708 337810 307760
rect 216490 306348 216496 306400
rect 216548 306388 216554 306400
rect 337654 306388 337660 306400
rect 216548 306360 337660 306388
rect 216548 306348 216554 306360
rect 337654 306348 337660 306360
rect 337712 306348 337718 306400
rect 321002 306280 321008 306332
rect 321060 306320 321066 306332
rect 337746 306320 337752 306332
rect 321060 306292 337752 306320
rect 321060 306280 321066 306292
rect 337746 306280 337752 306292
rect 337804 306280 337810 306332
rect 56502 304988 56508 305040
rect 56560 305028 56566 305040
rect 337654 305028 337660 305040
rect 56560 305000 337660 305028
rect 56560 304988 56566 305000
rect 337654 304988 337660 305000
rect 337712 304988 337718 305040
rect 169018 304920 169024 304972
rect 169076 304960 169082 304972
rect 337746 304960 337752 304972
rect 169076 304932 337752 304960
rect 169076 304920 169082 304932
rect 337746 304920 337752 304932
rect 337804 304920 337810 304972
rect 213822 303628 213828 303680
rect 213880 303668 213886 303680
rect 337654 303668 337660 303680
rect 213880 303640 337660 303668
rect 213880 303628 213886 303640
rect 337654 303628 337660 303640
rect 337712 303628 337718 303680
rect 333238 303560 333244 303612
rect 333296 303600 333302 303612
rect 336918 303600 336924 303612
rect 333296 303572 336924 303600
rect 333296 303560 333302 303572
rect 336918 303560 336924 303572
rect 336976 303560 336982 303612
rect 53742 302200 53748 302252
rect 53800 302240 53806 302252
rect 337654 302240 337660 302252
rect 53800 302212 337660 302240
rect 53800 302200 53806 302212
rect 337654 302200 337660 302212
rect 337712 302200 337718 302252
rect 166258 302132 166264 302184
rect 166316 302172 166322 302184
rect 337470 302172 337476 302184
rect 166316 302144 337476 302172
rect 166316 302132 166322 302144
rect 337470 302132 337476 302144
rect 337528 302132 337534 302184
rect 16850 301520 16856 301572
rect 16908 301560 16914 301572
rect 17126 301560 17132 301572
rect 16908 301532 17132 301560
rect 16908 301520 16914 301532
rect 17126 301520 17132 301532
rect 17184 301560 17190 301572
rect 17184 301532 26234 301560
rect 17184 301520 17190 301532
rect 26206 301492 26234 301532
rect 177206 301492 177212 301504
rect 26206 301464 177212 301492
rect 177206 301452 177212 301464
rect 177264 301452 177270 301504
rect 211062 300840 211068 300892
rect 211120 300880 211126 300892
rect 337654 300880 337660 300892
rect 211120 300852 337660 300880
rect 211120 300840 211126 300852
rect 337654 300840 337660 300852
rect 337712 300840 337718 300892
rect 327810 300772 327816 300824
rect 327868 300812 327874 300824
rect 337378 300812 337384 300824
rect 327868 300784 337384 300812
rect 327868 300772 327874 300784
rect 337378 300772 337384 300784
rect 337436 300772 337442 300824
rect 52362 299480 52368 299532
rect 52420 299520 52426 299532
rect 337654 299520 337660 299532
rect 52420 299492 337660 299520
rect 52420 299480 52426 299492
rect 337654 299480 337660 299492
rect 337712 299480 337718 299532
rect 162118 299412 162124 299464
rect 162176 299452 162182 299464
rect 337286 299452 337292 299464
rect 162176 299424 337292 299452
rect 162176 299412 162182 299424
rect 337286 299412 337292 299424
rect 337344 299412 337350 299464
rect 16758 298800 16764 298852
rect 16816 298840 16822 298852
rect 17218 298840 17224 298852
rect 16816 298812 17224 298840
rect 16816 298800 16822 298812
rect 17218 298800 17224 298812
rect 17276 298840 17282 298852
rect 17276 298812 26234 298840
rect 17276 298800 17282 298812
rect 26206 298772 26234 298812
rect 177390 298772 177396 298784
rect 26206 298744 177396 298772
rect 177390 298732 177396 298744
rect 177448 298732 177454 298784
rect 209314 298120 209320 298172
rect 209372 298160 209378 298172
rect 337102 298160 337108 298172
rect 209372 298132 337108 298160
rect 209372 298120 209378 298132
rect 337102 298120 337108 298132
rect 337160 298120 337166 298172
rect 200758 298052 200764 298104
rect 200816 298092 200822 298104
rect 336918 298092 336924 298104
rect 200816 298064 336924 298092
rect 200816 298052 200822 298064
rect 336918 298052 336924 298064
rect 336976 298052 336982 298104
rect 202138 297984 202144 298036
rect 202196 298024 202202 298036
rect 337654 298024 337660 298036
rect 202196 297996 337660 298024
rect 202196 297984 202202 297996
rect 337654 297984 337660 297996
rect 337712 297984 337718 298036
rect 178310 296828 178316 296880
rect 178368 296868 178374 296880
rect 197354 296868 197360 296880
rect 178368 296840 197360 296868
rect 178368 296828 178374 296840
rect 197354 296828 197360 296840
rect 197412 296828 197418 296880
rect 178402 296760 178408 296812
rect 178460 296800 178466 296812
rect 198734 296800 198740 296812
rect 178460 296772 198740 296800
rect 178460 296760 178466 296772
rect 198734 296760 198740 296772
rect 198792 296760 198798 296812
rect 48314 296692 48320 296744
rect 48372 296732 48378 296744
rect 337746 296732 337752 296744
rect 48372 296704 337752 296732
rect 48372 296692 48378 296704
rect 337746 296692 337752 296704
rect 337804 296692 337810 296744
rect 197354 296624 197360 296676
rect 197412 296664 197418 296676
rect 337102 296664 337108 296676
rect 197412 296636 337108 296664
rect 197412 296624 197418 296636
rect 337102 296624 337108 296636
rect 337160 296624 337166 296676
rect 198734 296556 198740 296608
rect 198792 296596 198798 296608
rect 337654 296596 337660 296608
rect 198792 296568 337660 296596
rect 198792 296556 198798 296568
rect 337654 296556 337660 296568
rect 337712 296556 337718 296608
rect 238018 295264 238024 295316
rect 238076 295304 238082 295316
rect 337654 295304 337660 295316
rect 238076 295276 337660 295304
rect 238076 295264 238082 295276
rect 337654 295264 337660 295276
rect 337712 295264 337718 295316
rect 239398 294652 239404 294704
rect 239456 294692 239462 294704
rect 316494 294692 316500 294704
rect 239456 294664 316500 294692
rect 239456 294652 239462 294664
rect 316494 294652 316500 294664
rect 316552 294652 316558 294704
rect 220630 294584 220636 294636
rect 220688 294624 220694 294636
rect 321002 294624 321008 294636
rect 220688 294596 321008 294624
rect 220688 294584 220694 294596
rect 321002 294584 321008 294596
rect 321060 294584 321066 294636
rect 178126 293972 178132 294024
rect 178184 294012 178190 294024
rect 204346 294012 204352 294024
rect 178184 293984 204352 294012
rect 178184 293972 178190 293984
rect 204346 293972 204352 293984
rect 204404 293972 204410 294024
rect 316494 293972 316500 294024
rect 316552 294012 316558 294024
rect 336918 294012 336924 294024
rect 316552 293984 336924 294012
rect 316552 293972 316558 293984
rect 336918 293972 336924 293984
rect 336976 293972 336982 294024
rect 3510 293904 3516 293956
rect 3568 293944 3574 293956
rect 327718 293944 327724 293956
rect 3568 293916 327724 293944
rect 3568 293904 3574 293916
rect 327718 293904 327724 293916
rect 327776 293904 327782 293956
rect 235258 293836 235264 293888
rect 235316 293876 235322 293888
rect 337746 293876 337752 293888
rect 235316 293848 337752 293876
rect 235316 293836 235322 293848
rect 337746 293836 337752 293848
rect 337804 293836 337810 293888
rect 236638 293768 236644 293820
rect 236696 293808 236702 293820
rect 337654 293808 337660 293820
rect 236696 293780 337660 293808
rect 236696 293768 236702 293780
rect 337654 293768 337660 293780
rect 337712 293768 337718 293820
rect 303062 293496 303068 293548
rect 303120 293536 303126 293548
rect 327810 293536 327816 293548
rect 303120 293508 327816 293536
rect 303120 293496 303126 293508
rect 327810 293496 327816 293508
rect 327868 293496 327874 293548
rect 266262 293428 266268 293480
rect 266320 293468 266326 293480
rect 325326 293468 325332 293480
rect 266320 293440 325332 293468
rect 266320 293428 266326 293440
rect 325326 293428 325332 293440
rect 325384 293428 325390 293480
rect 204346 293360 204352 293412
rect 204404 293400 204410 293412
rect 325142 293400 325148 293412
rect 204404 293372 325148 293400
rect 204404 293360 204410 293372
rect 325142 293360 325148 293372
rect 325200 293360 325206 293412
rect 213178 293292 213184 293344
rect 213236 293332 213242 293344
rect 336274 293332 336280 293344
rect 213236 293304 336280 293332
rect 213236 293292 213242 293304
rect 336274 293292 336280 293304
rect 336332 293292 336338 293344
rect 114462 293224 114468 293276
rect 114520 293264 114526 293276
rect 327994 293264 328000 293276
rect 114520 293236 328000 293264
rect 114520 293224 114526 293236
rect 327994 293224 328000 293236
rect 328052 293224 328058 293276
rect 234062 292476 234068 292528
rect 234120 292516 234126 292528
rect 337654 292516 337660 292528
rect 234120 292488 337660 292516
rect 234120 292476 234126 292488
rect 337654 292476 337660 292488
rect 337712 292476 337718 292528
rect 233878 292408 233884 292460
rect 233936 292448 233942 292460
rect 337746 292448 337752 292460
rect 233936 292420 337752 292448
rect 233936 292408 233942 292420
rect 337746 292408 337752 292420
rect 337804 292408 337810 292460
rect 262122 292340 262128 292392
rect 262180 292380 262186 292392
rect 323670 292380 323676 292392
rect 262180 292352 323676 292380
rect 262180 292340 262186 292352
rect 323670 292340 323676 292352
rect 323728 292340 323734 292392
rect 244182 292272 244188 292324
rect 244240 292312 244246 292324
rect 321278 292312 321284 292324
rect 244240 292284 321284 292312
rect 244240 292272 244246 292284
rect 321278 292272 321284 292284
rect 321336 292272 321342 292324
rect 237282 292204 237288 292256
rect 237340 292244 237346 292256
rect 322382 292244 322388 292256
rect 237340 292216 322388 292244
rect 237340 292204 237346 292216
rect 322382 292204 322388 292216
rect 322440 292204 322446 292256
rect 220446 292136 220452 292188
rect 220504 292176 220510 292188
rect 322474 292176 322480 292188
rect 220504 292148 322480 292176
rect 220504 292136 220510 292148
rect 322474 292136 322480 292148
rect 322532 292136 322538 292188
rect 216398 292068 216404 292120
rect 216456 292108 216462 292120
rect 332042 292108 332048 292120
rect 216456 292080 332048 292108
rect 216456 292068 216462 292080
rect 332042 292068 332048 292080
rect 332100 292068 332106 292120
rect 96522 292000 96528 292052
rect 96580 292040 96586 292052
rect 325510 292040 325516 292052
rect 96580 292012 325516 292040
rect 96580 292000 96586 292012
rect 325510 292000 325516 292012
rect 325568 292000 325574 292052
rect 78582 291932 78588 291984
rect 78640 291972 78646 291984
rect 332134 291972 332140 291984
rect 78640 291944 332140 291972
rect 78640 291932 78646 291944
rect 332134 291932 332140 291944
rect 332192 291932 332198 291984
rect 19794 291864 19800 291916
rect 19852 291904 19858 291916
rect 20070 291904 20076 291916
rect 19852 291876 20076 291904
rect 19852 291864 19858 291876
rect 20070 291864 20076 291876
rect 20128 291864 20134 291916
rect 73982 291864 73988 291916
rect 74040 291904 74046 291916
rect 329282 291904 329288 291916
rect 74040 291876 329288 291904
rect 74040 291864 74046 291876
rect 329282 291864 329288 291876
rect 329340 291864 329346 291916
rect 206278 291796 206284 291848
rect 206336 291836 206342 291848
rect 329190 291836 329196 291848
rect 206336 291808 329196 291836
rect 206336 291796 206342 291808
rect 329190 291796 329196 291808
rect 329248 291796 329254 291848
rect 284202 291728 284208 291780
rect 284260 291768 284266 291780
rect 330570 291768 330576 291780
rect 284260 291740 330576 291768
rect 284260 291728 284266 291740
rect 330570 291728 330576 291740
rect 330628 291728 330634 291780
rect 195974 291184 195980 291236
rect 196032 291224 196038 291236
rect 196158 291224 196164 291236
rect 196032 291196 196164 291224
rect 196032 291184 196038 291196
rect 196158 291184 196164 291196
rect 196216 291184 196222 291236
rect 106182 291116 106188 291168
rect 106240 291156 106246 291168
rect 336090 291156 336096 291168
rect 106240 291128 336096 291156
rect 106240 291116 106246 291128
rect 336090 291116 336096 291128
rect 336148 291116 336154 291168
rect 102042 291048 102048 291100
rect 102100 291088 102106 291100
rect 331858 291088 331864 291100
rect 102100 291060 331864 291088
rect 102100 291048 102106 291060
rect 331858 291048 331864 291060
rect 331916 291048 331922 291100
rect 104802 290980 104808 291032
rect 104860 291020 104866 291032
rect 334618 291020 334624 291032
rect 104860 290992 334624 291020
rect 104860 290980 104866 290992
rect 334618 290980 334624 290992
rect 334676 290980 334682 291032
rect 140682 290912 140688 290964
rect 140740 290952 140746 290964
rect 157518 290952 157524 290964
rect 140740 290924 157524 290952
rect 140740 290912 140746 290924
rect 157518 290912 157524 290924
rect 157576 290912 157582 290964
rect 316770 290912 316776 290964
rect 316828 290952 316834 290964
rect 337102 290952 337108 290964
rect 316828 290924 337108 290952
rect 316828 290912 316834 290924
rect 337102 290912 337108 290924
rect 337160 290912 337166 290964
rect 111702 290844 111708 290896
rect 111760 290884 111766 290896
rect 322290 290884 322296 290896
rect 111760 290856 322296 290884
rect 111760 290844 111766 290856
rect 322290 290844 322296 290856
rect 322348 290844 322354 290896
rect 118602 290776 118608 290828
rect 118660 290816 118666 290828
rect 318426 290816 318432 290828
rect 118660 290788 318432 290816
rect 118660 290776 118666 290788
rect 318426 290776 318432 290788
rect 318484 290776 318490 290828
rect 121362 290708 121368 290760
rect 121420 290748 121426 290760
rect 318334 290748 318340 290760
rect 121420 290720 318340 290748
rect 121420 290708 121426 290720
rect 318334 290708 318340 290720
rect 318392 290708 318398 290760
rect 122834 290640 122840 290692
rect 122892 290680 122898 290692
rect 318242 290680 318248 290692
rect 122892 290652 318248 290680
rect 122892 290640 122898 290652
rect 318242 290640 318248 290652
rect 318300 290640 318306 290692
rect 126882 290572 126888 290624
rect 126940 290612 126946 290624
rect 318150 290612 318156 290624
rect 126940 290584 318156 290612
rect 126940 290572 126946 290584
rect 318150 290572 318156 290584
rect 318208 290572 318214 290624
rect 139302 290504 139308 290556
rect 139360 290544 139366 290556
rect 157426 290544 157432 290556
rect 139360 290516 157432 290544
rect 139360 290504 139366 290516
rect 157426 290504 157432 290516
rect 157484 290504 157490 290556
rect 157518 290504 157524 290556
rect 157576 290544 157582 290556
rect 299658 290544 299664 290556
rect 157576 290516 299664 290544
rect 157576 290504 157582 290516
rect 299658 290504 299664 290516
rect 299716 290544 299722 290556
rect 317598 290544 317604 290556
rect 299716 290516 317604 290544
rect 299716 290504 299722 290516
rect 317598 290504 317604 290516
rect 317656 290544 317662 290556
rect 318610 290544 318616 290556
rect 317656 290516 318616 290544
rect 317656 290504 317662 290516
rect 318610 290504 318616 290516
rect 318668 290504 318674 290556
rect 151630 290436 151636 290488
rect 151688 290476 151694 290488
rect 160738 290476 160744 290488
rect 151688 290448 160744 290476
rect 151688 290436 151694 290448
rect 160738 290436 160744 290448
rect 160796 290476 160802 290488
rect 160796 290448 306374 290476
rect 160796 290436 160802 290448
rect 157426 290368 157432 290420
rect 157484 290408 157490 290420
rect 299014 290408 299020 290420
rect 157484 290380 299020 290408
rect 157484 290368 157490 290380
rect 299014 290368 299020 290380
rect 299072 290368 299078 290420
rect 306346 290408 306374 290448
rect 310790 290408 310796 290420
rect 306346 290380 310796 290408
rect 310790 290368 310796 290380
rect 310848 290408 310854 290420
rect 317414 290408 317420 290420
rect 310848 290380 317420 290408
rect 310848 290368 310854 290380
rect 317414 290368 317420 290380
rect 317472 290408 317478 290420
rect 318702 290408 318708 290420
rect 317472 290380 318708 290408
rect 317472 290368 317478 290380
rect 318702 290368 318708 290380
rect 318760 290368 318766 290420
rect 232498 290300 232504 290352
rect 232556 290340 232562 290352
rect 337470 290340 337476 290352
rect 232556 290312 337476 290340
rect 232556 290300 232562 290312
rect 337470 290300 337476 290312
rect 337528 290300 337534 290352
rect 234522 290232 234528 290284
rect 234580 290272 234586 290284
rect 318518 290272 318524 290284
rect 234580 290244 318524 290272
rect 234580 290232 234586 290244
rect 318518 290232 318524 290244
rect 318576 290232 318582 290284
rect 286594 290164 286600 290216
rect 286652 290204 286658 290216
rect 319438 290204 319444 290216
rect 286652 290176 319444 290204
rect 286652 290164 286658 290176
rect 319438 290164 319444 290176
rect 319496 290164 319502 290216
rect 108942 290096 108948 290148
rect 109000 290136 109006 290148
rect 320910 290136 320916 290148
rect 109000 290108 320916 290136
rect 109000 290096 109006 290108
rect 320910 290096 320916 290108
rect 320968 290096 320974 290148
rect 178126 289824 178132 289876
rect 178184 289864 178190 289876
rect 204254 289864 204260 289876
rect 178184 289836 204260 289864
rect 178184 289824 178190 289836
rect 204254 289824 204260 289836
rect 204312 289864 204318 289876
rect 204714 289864 204720 289876
rect 204312 289836 204720 289864
rect 204312 289824 204318 289836
rect 204714 289824 204720 289836
rect 204772 289824 204778 289876
rect 229002 289756 229008 289808
rect 229060 289796 229066 289808
rect 337746 289796 337752 289808
rect 229060 289768 337752 289796
rect 229060 289756 229066 289768
rect 337746 289756 337752 289768
rect 337804 289756 337810 289808
rect 229738 289688 229744 289740
rect 229796 289728 229802 289740
rect 337654 289728 337660 289740
rect 229796 289700 337660 289728
rect 229796 289688 229802 289700
rect 337654 289688 337660 289700
rect 337712 289688 337718 289740
rect 299014 289620 299020 289672
rect 299072 289660 299078 289672
rect 317506 289660 317512 289672
rect 299072 289632 317512 289660
rect 299072 289620 299078 289632
rect 317506 289620 317512 289632
rect 317564 289660 317570 289672
rect 327718 289660 327724 289672
rect 317564 289632 327724 289660
rect 317564 289620 317570 289632
rect 327718 289620 327724 289632
rect 327776 289620 327782 289672
rect 302878 289552 302884 289604
rect 302936 289592 302942 289604
rect 318150 289592 318156 289604
rect 302936 289564 318156 289592
rect 302936 289552 302942 289564
rect 318150 289552 318156 289564
rect 318208 289552 318214 289604
rect 222838 289484 222844 289536
rect 222896 289524 222902 289536
rect 317414 289524 317420 289536
rect 222896 289496 317420 289524
rect 222896 289484 222902 289496
rect 317414 289484 317420 289496
rect 317472 289484 317478 289536
rect 215110 289416 215116 289468
rect 215168 289456 215174 289468
rect 322014 289456 322020 289468
rect 215168 289428 322020 289456
rect 215168 289416 215174 289428
rect 322014 289416 322020 289428
rect 322072 289416 322078 289468
rect 16666 289348 16672 289400
rect 16724 289388 16730 289400
rect 70394 289388 70400 289400
rect 16724 289360 70400 289388
rect 16724 289348 16730 289360
rect 70394 289348 70400 289360
rect 70452 289348 70458 289400
rect 217870 289348 217876 289400
rect 217928 289388 217934 289400
rect 324314 289388 324320 289400
rect 217928 289360 324320 289388
rect 217928 289348 217934 289360
rect 324314 289348 324320 289360
rect 324372 289348 324378 289400
rect 17954 289280 17960 289332
rect 18012 289320 18018 289332
rect 74534 289320 74540 289332
rect 18012 289292 74540 289320
rect 18012 289280 18018 289292
rect 74534 289280 74540 289292
rect 74592 289280 74598 289332
rect 204714 289280 204720 289332
rect 204772 289320 204778 289332
rect 331858 289320 331864 289332
rect 204772 289292 331864 289320
rect 204772 289280 204778 289292
rect 331858 289280 331864 289292
rect 331916 289280 331922 289332
rect 17218 289212 17224 289264
rect 17276 289252 17282 289264
rect 77294 289252 77300 289264
rect 17276 289224 77300 289252
rect 17276 289212 17282 289224
rect 77294 289212 77300 289224
rect 77352 289212 77358 289264
rect 177114 289212 177120 289264
rect 177172 289252 177178 289264
rect 337470 289252 337476 289264
rect 177172 289224 337476 289252
rect 177172 289212 177178 289224
rect 337470 289212 337476 289224
rect 337528 289212 337534 289264
rect 17034 289144 17040 289196
rect 17092 289184 17098 289196
rect 336734 289184 336740 289196
rect 17092 289156 336740 289184
rect 17092 289144 17098 289156
rect 336734 289144 336740 289156
rect 336792 289144 336798 289196
rect 17126 289076 17132 289128
rect 17184 289116 17190 289128
rect 78674 289116 78680 289128
rect 17184 289088 78680 289116
rect 17184 289076 17190 289088
rect 78674 289076 78680 289088
rect 78732 289076 78738 289128
rect 318702 289076 318708 289128
rect 318760 289116 318766 289128
rect 338758 289116 338764 289128
rect 318760 289088 338764 289116
rect 318760 289076 318766 289088
rect 338758 289076 338764 289088
rect 338816 289076 338822 289128
rect 180702 289008 180708 289060
rect 180760 289048 180766 289060
rect 195974 289048 195980 289060
rect 180760 289020 195980 289048
rect 180760 289008 180766 289020
rect 195974 289008 195980 289020
rect 196032 289008 196038 289060
rect 178034 288940 178040 288992
rect 178092 288980 178098 288992
rect 196066 288980 196072 288992
rect 178092 288952 196072 288980
rect 178092 288940 178098 288952
rect 196066 288940 196072 288952
rect 196124 288940 196130 288992
rect 177482 288872 177488 288924
rect 177540 288912 177546 288924
rect 337562 288912 337568 288924
rect 177540 288884 337568 288912
rect 177540 288872 177546 288884
rect 337562 288872 337568 288884
rect 337620 288872 337626 288924
rect 177206 288804 177212 288856
rect 177264 288844 177270 288856
rect 337378 288844 337384 288856
rect 177264 288816 337384 288844
rect 177264 288804 177270 288816
rect 337378 288804 337384 288816
rect 337436 288804 337442 288856
rect 177574 288736 177580 288788
rect 177632 288776 177638 288788
rect 337841 288779 337899 288785
rect 337841 288776 337853 288779
rect 177632 288748 337853 288776
rect 177632 288736 177638 288748
rect 337841 288745 337853 288748
rect 337887 288745 337899 288779
rect 337841 288739 337899 288745
rect 177666 288668 177672 288720
rect 177724 288708 177730 288720
rect 338022 288708 338028 288720
rect 177724 288680 338028 288708
rect 177724 288668 177730 288680
rect 338022 288668 338028 288680
rect 338080 288668 338086 288720
rect 177114 288600 177120 288652
rect 177172 288640 177178 288652
rect 177482 288640 177488 288652
rect 177172 288612 177488 288640
rect 177172 288600 177178 288612
rect 177482 288600 177488 288612
rect 177540 288600 177546 288652
rect 177758 288600 177764 288652
rect 177816 288640 177822 288652
rect 337930 288640 337936 288652
rect 177816 288612 337936 288640
rect 177816 288600 177822 288612
rect 337930 288600 337936 288612
rect 337988 288600 337994 288652
rect 177298 288532 177304 288584
rect 177356 288572 177362 288584
rect 337838 288572 337844 288584
rect 177356 288544 337844 288572
rect 177356 288532 177362 288544
rect 337838 288532 337844 288544
rect 337896 288532 337902 288584
rect 177482 288464 177488 288516
rect 177540 288504 177546 288516
rect 177758 288504 177764 288516
rect 177540 288476 177764 288504
rect 177540 288464 177546 288476
rect 177758 288464 177764 288476
rect 177816 288464 177822 288516
rect 177850 288464 177856 288516
rect 177908 288504 177914 288516
rect 336826 288504 336832 288516
rect 177908 288476 336832 288504
rect 177908 288464 177914 288476
rect 336826 288464 336832 288476
rect 336884 288464 336890 288516
rect 160002 288396 160008 288448
rect 160060 288436 160066 288448
rect 320910 288436 320916 288448
rect 160060 288408 320916 288436
rect 160060 288396 160066 288408
rect 320910 288396 320916 288408
rect 320968 288396 320974 288448
rect 225598 288328 225604 288380
rect 225656 288368 225662 288380
rect 336918 288368 336924 288380
rect 225656 288340 336924 288368
rect 225656 288328 225662 288340
rect 336918 288328 336924 288340
rect 336976 288328 336982 288380
rect 226978 288260 226984 288312
rect 227036 288300 227042 288312
rect 337654 288300 337660 288312
rect 227036 288272 337660 288300
rect 227036 288260 227042 288272
rect 337654 288260 337660 288272
rect 337712 288260 337718 288312
rect 227530 288192 227536 288244
rect 227588 288232 227594 288244
rect 337746 288232 337752 288244
rect 227588 288204 337752 288232
rect 227588 288192 227594 288204
rect 337746 288192 337752 288204
rect 337804 288192 337810 288244
rect 211982 287988 211988 288040
rect 212040 288028 212046 288040
rect 337194 288028 337200 288040
rect 212040 288000 337200 288028
rect 212040 287988 212046 288000
rect 337194 287988 337200 288000
rect 337252 287988 337258 288040
rect 211798 287920 211804 287972
rect 211856 287960 211862 287972
rect 337286 287960 337292 287972
rect 211856 287932 337292 287960
rect 211856 287920 211862 287932
rect 337286 287920 337292 287932
rect 337344 287920 337350 287972
rect 19337 287895 19395 287901
rect 19337 287861 19349 287895
rect 19383 287892 19395 287895
rect 36538 287892 36544 287904
rect 19383 287864 36544 287892
rect 19383 287861 19395 287864
rect 19337 287855 19395 287861
rect 36538 287852 36544 287864
rect 36596 287852 36602 287904
rect 209038 287852 209044 287904
rect 209096 287892 209102 287904
rect 334618 287892 334624 287904
rect 209096 287864 334624 287892
rect 209096 287852 209102 287864
rect 334618 287852 334624 287864
rect 334676 287852 334682 287904
rect 19426 287784 19432 287836
rect 19484 287824 19490 287836
rect 37918 287824 37924 287836
rect 19484 287796 37924 287824
rect 19484 287784 19490 287796
rect 37918 287784 37924 287796
rect 37976 287784 37982 287836
rect 210418 287784 210424 287836
rect 210476 287824 210482 287836
rect 337102 287824 337108 287836
rect 210476 287796 337108 287824
rect 210476 287784 210482 287796
rect 337102 287784 337108 287796
rect 337160 287784 337166 287836
rect 19334 287716 19340 287768
rect 19392 287756 19398 287768
rect 40678 287756 40684 287768
rect 19392 287728 40684 287756
rect 19392 287716 19398 287728
rect 40678 287716 40684 287728
rect 40736 287716 40742 287768
rect 195974 287716 195980 287768
rect 196032 287756 196038 287768
rect 337010 287756 337016 287768
rect 196032 287728 337016 287756
rect 196032 287716 196038 287728
rect 337010 287716 337016 287728
rect 337068 287716 337074 287768
rect 18046 287648 18052 287700
rect 18104 287688 18110 287700
rect 42058 287688 42064 287700
rect 18104 287660 42064 287688
rect 18104 287648 18110 287660
rect 42058 287648 42064 287660
rect 42116 287648 42122 287700
rect 196066 287648 196072 287700
rect 196124 287688 196130 287700
rect 337562 287688 337568 287700
rect 196124 287660 337568 287688
rect 196124 287648 196130 287660
rect 337562 287648 337568 287660
rect 337620 287648 337626 287700
rect 336734 287580 336740 287632
rect 336792 287620 336798 287632
rect 337654 287620 337660 287632
rect 336792 287592 337660 287620
rect 336792 287580 336798 287592
rect 337654 287580 337660 287592
rect 337712 287580 337718 287632
rect 178773 287419 178831 287425
rect 142126 287388 151814 287416
rect 16942 287308 16948 287360
rect 17000 287348 17006 287360
rect 142126 287348 142154 287388
rect 17000 287320 142154 287348
rect 17000 287308 17006 287320
rect 150894 287308 150900 287360
rect 150952 287348 150958 287360
rect 151630 287348 151636 287360
rect 150952 287320 151636 287348
rect 150952 287308 150958 287320
rect 151630 287308 151636 287320
rect 151688 287308 151694 287360
rect 151786 287348 151814 287388
rect 178773 287385 178785 287419
rect 178819 287416 178831 287419
rect 180334 287416 180340 287428
rect 178819 287388 180340 287416
rect 178819 287385 178831 287388
rect 178773 287379 178831 287385
rect 180334 287376 180340 287388
rect 180392 287376 180398 287428
rect 180702 287416 180708 287428
rect 180663 287388 180708 287416
rect 180702 287376 180708 287388
rect 180760 287376 180766 287428
rect 318058 287348 318064 287360
rect 151786 287320 318064 287348
rect 318058 287308 318064 287320
rect 318116 287308 318122 287360
rect 151648 287280 151676 287308
rect 157978 287280 157984 287292
rect 151648 287252 157984 287280
rect 157978 287240 157984 287252
rect 158036 287240 158042 287292
rect 177850 287240 177856 287292
rect 177908 287280 177914 287292
rect 322290 287280 322296 287292
rect 177908 287252 322296 287280
rect 177908 287240 177914 287252
rect 322290 287240 322296 287252
rect 322348 287240 322354 287292
rect 337930 287280 337936 287292
rect 337891 287252 337936 287280
rect 337930 287240 337936 287252
rect 337988 287240 337994 287292
rect 338022 287240 338028 287292
rect 338080 287240 338086 287292
rect 338040 287088 338068 287240
rect 337841 287079 337899 287085
rect 337841 287045 337853 287079
rect 337887 287076 337899 287079
rect 337930 287076 337936 287088
rect 337887 287048 337936 287076
rect 337887 287045 337899 287048
rect 337841 287039 337899 287045
rect 337930 287036 337936 287048
rect 337988 287036 337994 287088
rect 338022 287036 338028 287088
rect 338080 287036 338086 287088
rect 19426 286968 19432 287020
rect 19484 287008 19490 287020
rect 19981 287011 20039 287017
rect 19981 287008 19993 287011
rect 19484 286980 19993 287008
rect 19484 286968 19490 286980
rect 19981 286977 19993 286980
rect 20027 286977 20039 287011
rect 19981 286971 20039 286977
rect 316678 286968 316684 287020
rect 316736 287008 316742 287020
rect 337194 287008 337200 287020
rect 316736 286980 336780 287008
rect 316736 286968 316742 286980
rect 336752 286952 336780 286980
rect 336844 286980 337200 287008
rect 317414 286900 317420 286952
rect 317472 286940 317478 286952
rect 317472 286912 335354 286940
rect 317472 286900 317478 286912
rect 19334 286804 19340 286816
rect 19295 286776 19340 286804
rect 19334 286764 19340 286776
rect 19392 286764 19398 286816
rect 335326 286804 335354 286912
rect 336734 286900 336740 286952
rect 336792 286900 336798 286952
rect 336844 286884 336872 286980
rect 337194 286968 337200 286980
rect 337252 286968 337258 287020
rect 336826 286832 336832 286884
rect 336884 286832 336890 286884
rect 337102 286872 337108 286884
rect 337063 286844 337108 286872
rect 337102 286832 337108 286844
rect 337160 286832 337166 286884
rect 337194 286832 337200 286884
rect 337252 286872 337258 286884
rect 338114 286872 338120 286884
rect 337252 286844 338120 286872
rect 337252 286832 337258 286844
rect 338114 286832 338120 286844
rect 338172 286832 338178 286884
rect 337470 286804 337476 286816
rect 335326 286776 337476 286804
rect 337470 286764 337476 286776
rect 337528 286764 337534 286816
rect 337930 286804 337936 286816
rect 337891 286776 337936 286804
rect 337930 286764 337936 286776
rect 337988 286764 337994 286816
rect 337010 285744 337016 285796
rect 337068 285784 337074 285796
rect 337654 285784 337660 285796
rect 337068 285756 337660 285784
rect 337068 285744 337074 285756
rect 337654 285744 337660 285756
rect 337712 285744 337718 285796
rect 336734 285676 336740 285728
rect 336792 285716 336798 285728
rect 337286 285716 337292 285728
rect 336792 285688 337292 285716
rect 336792 285676 336798 285688
rect 337286 285676 337292 285688
rect 337344 285676 337350 285728
rect 322474 285608 322480 285660
rect 322532 285648 322538 285660
rect 337654 285648 337660 285660
rect 322532 285620 337660 285648
rect 322532 285608 322538 285620
rect 337654 285608 337660 285620
rect 337712 285608 337718 285660
rect 323854 285540 323860 285592
rect 323912 285580 323918 285592
rect 337286 285580 337292 285592
rect 323912 285552 337292 285580
rect 323912 285540 323918 285552
rect 337286 285540 337292 285552
rect 337344 285540 337350 285592
rect 336642 285132 336648 285184
rect 336700 285172 336706 285184
rect 337286 285172 337292 285184
rect 336700 285144 337292 285172
rect 336700 285132 336706 285144
rect 337286 285132 337292 285144
rect 337344 285132 337350 285184
rect 337470 284316 337476 284368
rect 337528 284356 337534 284368
rect 337746 284356 337752 284368
rect 337528 284328 337752 284356
rect 337528 284316 337534 284328
rect 337746 284316 337752 284328
rect 337804 284316 337810 284368
rect 321002 284248 321008 284300
rect 321060 284288 321066 284300
rect 337654 284288 337660 284300
rect 321060 284260 337660 284288
rect 321060 284248 321066 284260
rect 337654 284248 337660 284260
rect 337712 284248 337718 284300
rect 327902 284180 327908 284232
rect 327960 284220 327966 284232
rect 337746 284220 337752 284232
rect 327960 284192 337752 284220
rect 327960 284180 327966 284192
rect 337746 284180 337752 284192
rect 337804 284180 337810 284232
rect 178678 283064 178684 283076
rect 178639 283036 178684 283064
rect 178678 283024 178684 283036
rect 178736 283024 178742 283076
rect 178678 282888 178684 282940
rect 178736 282928 178742 282940
rect 178773 282931 178831 282937
rect 178773 282928 178785 282931
rect 178736 282900 178785 282928
rect 178736 282888 178742 282900
rect 178773 282897 178785 282900
rect 178819 282897 178831 282931
rect 178773 282891 178831 282897
rect 324314 282820 324320 282872
rect 324372 282860 324378 282872
rect 337654 282860 337660 282872
rect 324372 282832 337660 282860
rect 324372 282820 324378 282832
rect 337654 282820 337660 282832
rect 337712 282820 337718 282872
rect 332042 282752 332048 282804
rect 332100 282792 332106 282804
rect 337746 282792 337752 282804
rect 332100 282764 337752 282792
rect 332100 282752 332106 282764
rect 337746 282752 337752 282764
rect 337804 282752 337810 282804
rect 337105 282591 337163 282597
rect 337105 282557 337117 282591
rect 337151 282588 337163 282591
rect 337654 282588 337660 282600
rect 337151 282560 337660 282588
rect 337151 282557 337163 282560
rect 337105 282551 337163 282557
rect 337654 282548 337660 282560
rect 337712 282548 337718 282600
rect 337286 282344 337292 282396
rect 337344 282384 337350 282396
rect 337344 282356 337424 282384
rect 337344 282344 337350 282356
rect 337396 282192 337424 282356
rect 337378 282140 337384 282192
rect 337436 282140 337442 282192
rect 322014 281392 322020 281444
rect 322072 281432 322078 281444
rect 337654 281432 337660 281444
rect 322072 281404 337660 281432
rect 322072 281392 322078 281404
rect 337654 281392 337660 281404
rect 337712 281392 337718 281444
rect 334618 278672 334624 278724
rect 334676 278712 334682 278724
rect 337654 278712 337660 278724
rect 334676 278684 337660 278712
rect 334676 278672 334682 278684
rect 337654 278672 337660 278684
rect 337712 278672 337718 278724
rect 330662 278604 330668 278656
rect 330720 278644 330726 278656
rect 337746 278644 337752 278656
rect 330720 278616 337752 278644
rect 330720 278604 330726 278616
rect 337746 278604 337752 278616
rect 337804 278604 337810 278656
rect 337654 278060 337660 278112
rect 337712 278100 337718 278112
rect 338022 278100 338028 278112
rect 337712 278072 338028 278100
rect 337712 278060 337718 278072
rect 338022 278060 338028 278072
rect 338080 278060 338086 278112
rect 337378 277924 337384 277976
rect 337436 277964 337442 277976
rect 338022 277964 338028 277976
rect 337436 277936 338028 277964
rect 337436 277924 337442 277936
rect 338022 277924 338028 277936
rect 338080 277924 338086 277976
rect 337102 277584 337108 277636
rect 337160 277584 337166 277636
rect 337194 277584 337200 277636
rect 337252 277624 337258 277636
rect 337252 277596 337792 277624
rect 337252 277584 337258 277596
rect 19426 277488 19432 277500
rect 19387 277460 19432 277488
rect 19426 277448 19432 277460
rect 19484 277448 19490 277500
rect 337120 277432 337148 277584
rect 337764 277432 337792 277596
rect 337102 277380 337108 277432
rect 337160 277380 337166 277432
rect 337746 277380 337752 277432
rect 337804 277380 337810 277432
rect 19426 277352 19432 277364
rect 19387 277324 19432 277352
rect 19426 277312 19432 277324
rect 19484 277312 19490 277364
rect 331858 277312 331864 277364
rect 331916 277352 331922 277364
rect 337378 277352 337384 277364
rect 331916 277324 337384 277352
rect 331916 277312 331922 277324
rect 337378 277312 337384 277324
rect 337436 277312 337442 277364
rect 329190 277244 329196 277296
rect 329248 277284 329254 277296
rect 337838 277284 337844 277296
rect 329248 277256 337844 277284
rect 329248 277244 329254 277256
rect 337838 277244 337844 277256
rect 337896 277244 337902 277296
rect 325142 275952 325148 276004
rect 325200 275992 325206 276004
rect 337838 275992 337844 276004
rect 325200 275964 337844 275992
rect 325200 275952 325206 275964
rect 337838 275952 337844 275964
rect 337896 275952 337902 276004
rect 334802 275884 334808 275936
rect 334860 275924 334866 275936
rect 337378 275924 337384 275936
rect 334860 275896 337384 275924
rect 334860 275884 334866 275896
rect 337378 275884 337384 275896
rect 337436 275884 337442 275936
rect 322290 274592 322296 274644
rect 322348 274632 322354 274644
rect 337838 274632 337844 274644
rect 322348 274604 337844 274632
rect 322348 274592 322354 274604
rect 337838 274592 337844 274604
rect 337896 274592 337902 274644
rect 482370 273776 482376 273828
rect 482428 273816 482434 273828
rect 485038 273816 485044 273828
rect 482428 273788 485044 273816
rect 482428 273776 482434 273788
rect 485038 273776 485044 273788
rect 485096 273776 485102 273828
rect 318058 273164 318064 273216
rect 318116 273204 318122 273216
rect 337838 273204 337844 273216
rect 318116 273176 337844 273204
rect 318116 273164 318122 273176
rect 337838 273164 337844 273176
rect 337896 273164 337902 273216
rect 482278 273164 482284 273216
rect 482336 273204 482342 273216
rect 580166 273204 580172 273216
rect 482336 273176 580172 273204
rect 482336 273164 482342 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 319438 271804 319444 271856
rect 319496 271844 319502 271856
rect 337838 271844 337844 271856
rect 319496 271816 337844 271844
rect 319496 271804 319502 271816
rect 337838 271804 337844 271816
rect 337896 271804 337902 271856
rect 323762 271736 323768 271788
rect 323820 271776 323826 271788
rect 337102 271776 337108 271788
rect 323820 271748 337108 271776
rect 323820 271736 323826 271748
rect 337102 271736 337108 271748
rect 337160 271736 337166 271788
rect 320910 270376 320916 270428
rect 320968 270416 320974 270428
rect 337838 270416 337844 270428
rect 320968 270388 337844 270416
rect 320968 270376 320974 270388
rect 337838 270376 337844 270388
rect 337896 270376 337902 270428
rect 178678 267628 178684 267640
rect 178639 267600 178684 267628
rect 178678 267588 178684 267600
rect 178736 267588 178742 267640
rect 481910 264936 481916 264988
rect 481968 264976 481974 264988
rect 483658 264976 483664 264988
rect 481968 264948 483664 264976
rect 481968 264936 481974 264948
rect 483658 264936 483664 264948
rect 483716 264936 483722 264988
rect 327810 262896 327816 262948
rect 327868 262936 327874 262948
rect 336826 262936 336832 262948
rect 327868 262908 336832 262936
rect 327868 262896 327874 262908
rect 336826 262896 336832 262908
rect 336884 262936 336890 262948
rect 337378 262936 337384 262948
rect 336884 262908 337384 262936
rect 336884 262896 336890 262908
rect 337378 262896 337384 262908
rect 337436 262896 337442 262948
rect 318150 262828 318156 262880
rect 318208 262868 318214 262880
rect 337010 262868 337016 262880
rect 318208 262840 337016 262868
rect 318208 262828 318214 262840
rect 337010 262828 337016 262840
rect 337068 262868 337074 262880
rect 337470 262868 337476 262880
rect 337068 262840 337476 262868
rect 337068 262828 337074 262840
rect 337470 262828 337476 262840
rect 337528 262828 337534 262880
rect 319438 262148 319444 262200
rect 319496 262188 319502 262200
rect 319898 262188 319904 262200
rect 319496 262160 319904 262188
rect 319496 262148 319502 262160
rect 319898 262148 319904 262160
rect 319956 262148 319962 262200
rect 319806 261536 319812 261588
rect 319864 261576 319870 261588
rect 337654 261576 337660 261588
rect 319864 261548 337660 261576
rect 319864 261536 319870 261548
rect 337654 261536 337660 261548
rect 337712 261536 337718 261588
rect 319438 261468 319444 261520
rect 319496 261508 319502 261520
rect 337470 261508 337476 261520
rect 319496 261480 337476 261508
rect 319496 261468 319502 261480
rect 337470 261468 337476 261480
rect 337528 261468 337534 261520
rect 319530 260244 319536 260296
rect 319588 260284 319594 260296
rect 337102 260284 337108 260296
rect 319588 260256 337108 260284
rect 319588 260244 319594 260256
rect 337102 260244 337108 260256
rect 337160 260244 337166 260296
rect 319714 260176 319720 260228
rect 319772 260216 319778 260228
rect 337746 260216 337752 260228
rect 319772 260188 337752 260216
rect 319772 260176 319778 260188
rect 337746 260176 337752 260188
rect 337804 260176 337810 260228
rect 319622 260108 319628 260160
rect 319680 260148 319686 260160
rect 337654 260148 337660 260160
rect 319680 260120 337660 260148
rect 319680 260108 319686 260120
rect 337654 260108 337660 260120
rect 337712 260108 337718 260160
rect 318610 259360 318616 259412
rect 318668 259400 318674 259412
rect 337654 259400 337660 259412
rect 318668 259372 337660 259400
rect 318668 259360 318674 259372
rect 337654 259360 337660 259372
rect 337712 259360 337718 259412
rect 482002 259360 482008 259412
rect 482060 259400 482066 259412
rect 580166 259400 580172 259412
rect 482060 259372 580172 259400
rect 482060 259360 482066 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 327718 259292 327724 259344
rect 327776 259332 327782 259344
rect 336918 259332 336924 259344
rect 327776 259304 336924 259332
rect 327776 259292 327782 259304
rect 336918 259292 336924 259304
rect 336976 259292 336982 259344
rect 338758 258204 338764 258256
rect 338816 258244 338822 258256
rect 340322 258244 340328 258256
rect 338816 258216 340328 258244
rect 338816 258204 338822 258216
rect 340322 258204 340328 258216
rect 340380 258204 340386 258256
rect 19426 258176 19432 258188
rect 19387 258148 19432 258176
rect 19426 258136 19432 258148
rect 19484 258136 19490 258188
rect 178678 258108 178684 258120
rect 178639 258080 178684 258108
rect 178678 258068 178684 258080
rect 178736 258068 178742 258120
rect 179598 258074 179604 258086
rect 19426 258040 19432 258052
rect 19387 258012 19432 258040
rect 19426 258000 19432 258012
rect 19484 258000 19490 258052
rect 179545 258046 179604 258074
rect 179598 258034 179604 258046
rect 179656 258034 179662 258086
rect 179601 258009 179613 258034
rect 179647 258009 179659 258034
rect 179601 258003 179659 258009
rect 336918 258000 336924 258052
rect 336976 258040 336982 258052
rect 339034 258040 339040 258052
rect 336976 258012 339040 258040
rect 336976 258000 336982 258012
rect 339034 258000 339040 258012
rect 339092 258000 339098 258052
rect 178678 257972 178684 257984
rect 178639 257944 178684 257972
rect 178678 257932 178684 257944
rect 178736 257932 178742 257984
rect 179690 257796 179696 257848
rect 179748 257836 179754 257848
rect 179969 257839 180027 257845
rect 179969 257836 179981 257839
rect 179748 257808 179981 257836
rect 179748 257796 179754 257808
rect 179969 257805 179981 257808
rect 180015 257805 180027 257839
rect 179969 257799 180027 257805
rect 336090 256572 336096 256624
rect 336148 256612 336154 256624
rect 345934 256612 345940 256624
rect 336148 256584 345940 256612
rect 336148 256572 336154 256584
rect 345934 256572 345940 256584
rect 345992 256572 345998 256624
rect 347038 256572 347044 256624
rect 347096 256612 347102 256624
rect 365714 256612 365720 256624
rect 347096 256584 365720 256612
rect 347096 256572 347102 256584
rect 365714 256572 365720 256584
rect 365772 256572 365778 256624
rect 327718 256504 327724 256556
rect 327776 256544 327782 256556
rect 361574 256544 361580 256556
rect 327776 256516 361580 256544
rect 327776 256504 327782 256516
rect 361574 256504 361580 256516
rect 361632 256504 361638 256556
rect 331858 256436 331864 256488
rect 331916 256476 331922 256488
rect 367094 256476 367100 256488
rect 331916 256448 367100 256476
rect 331916 256436 331922 256448
rect 367094 256436 367100 256448
rect 367152 256436 367158 256488
rect 367738 256436 367744 256488
rect 367796 256476 367802 256488
rect 369302 256476 369308 256488
rect 367796 256448 369308 256476
rect 367796 256436 367802 256448
rect 369302 256436 369308 256448
rect 369360 256436 369366 256488
rect 374638 256436 374644 256488
rect 374696 256476 374702 256488
rect 390554 256476 390560 256488
rect 374696 256448 390560 256476
rect 374696 256436 374702 256448
rect 390554 256436 390560 256448
rect 390612 256436 390618 256488
rect 334618 256368 334624 256420
rect 334676 256408 334682 256420
rect 379882 256408 379888 256420
rect 334676 256380 379888 256408
rect 334676 256368 334682 256380
rect 379882 256368 379888 256380
rect 379940 256368 379946 256420
rect 320910 256300 320916 256352
rect 320968 256340 320974 256352
rect 350810 256340 350816 256352
rect 320968 256312 350816 256340
rect 320968 256300 320974 256312
rect 350810 256300 350816 256312
rect 350868 256300 350874 256352
rect 352558 256300 352564 256352
rect 352616 256340 352622 256352
rect 408954 256340 408960 256352
rect 352616 256312 408960 256340
rect 352616 256300 352622 256312
rect 408954 256300 408960 256312
rect 409012 256300 409018 256352
rect 475378 256300 475384 256352
rect 475436 256340 475442 256352
rect 477678 256340 477684 256352
rect 475436 256312 477684 256340
rect 475436 256300 475442 256312
rect 477678 256300 477684 256312
rect 477736 256300 477742 256352
rect 340230 256232 340236 256284
rect 340288 256272 340294 256284
rect 397454 256272 397460 256284
rect 340288 256244 397460 256272
rect 340288 256232 340294 256244
rect 397454 256232 397460 256244
rect 397512 256232 397518 256284
rect 318058 256164 318064 256216
rect 318116 256204 318122 256216
rect 404998 256204 405004 256216
rect 318116 256176 405004 256204
rect 318116 256164 318122 256176
rect 404998 256164 405004 256176
rect 405056 256164 405062 256216
rect 322290 256096 322296 256148
rect 322348 256136 322354 256148
rect 415578 256136 415584 256148
rect 322348 256108 415584 256136
rect 322348 256096 322354 256108
rect 415578 256096 415584 256108
rect 415636 256096 415642 256148
rect 436738 256096 436744 256148
rect 436796 256136 436802 256148
rect 473722 256136 473728 256148
rect 436796 256108 473728 256136
rect 436796 256096 436802 256108
rect 473722 256096 473728 256108
rect 473780 256096 473786 256148
rect 323670 256028 323676 256080
rect 323728 256068 323734 256080
rect 455414 256068 455420 256080
rect 323728 256040 455420 256068
rect 323728 256028 323734 256040
rect 455414 256028 455420 256040
rect 455472 256028 455478 256080
rect 324958 255960 324964 256012
rect 325016 256000 325022 256012
rect 463142 256000 463148 256012
rect 325016 255972 463148 256000
rect 325016 255960 325022 255972
rect 463142 255960 463148 255972
rect 463200 255960 463206 256012
rect 465718 255960 465724 256012
rect 465776 256000 465782 256012
rect 475010 256000 475016 256012
rect 465776 255972 475016 256000
rect 465776 255960 465782 255972
rect 475010 255960 475016 255972
rect 475068 255960 475074 256012
rect 340138 255892 340144 255944
rect 340196 255932 340202 255944
rect 344278 255932 344284 255944
rect 340196 255904 344284 255932
rect 340196 255892 340202 255904
rect 344278 255892 344284 255904
rect 344336 255892 344342 255944
rect 339402 255756 339408 255808
rect 339460 255796 339466 255808
rect 340874 255796 340880 255808
rect 339460 255768 340880 255796
rect 339460 255756 339466 255768
rect 340874 255756 340880 255768
rect 340932 255796 340938 255808
rect 341610 255796 341616 255808
rect 340932 255768 341616 255796
rect 340932 255756 340938 255768
rect 341610 255756 341616 255768
rect 341668 255756 341674 255808
rect 370498 255620 370504 255672
rect 370556 255660 370562 255672
rect 373258 255660 373264 255672
rect 370556 255632 373264 255660
rect 370556 255620 370562 255632
rect 373258 255620 373264 255632
rect 373316 255620 373322 255672
rect 345658 255484 345664 255536
rect 345716 255524 345722 255536
rect 348234 255524 348240 255536
rect 345716 255496 348240 255524
rect 345716 255484 345722 255496
rect 348234 255484 348240 255496
rect 348292 255484 348298 255536
rect 338850 255348 338856 255400
rect 338908 255388 338914 255400
rect 346854 255388 346860 255400
rect 338908 255360 346860 255388
rect 338908 255348 338914 255360
rect 346854 255348 346860 255360
rect 346912 255348 346918 255400
rect 179690 253852 179696 253904
rect 179748 253892 179754 253904
rect 179969 253895 180027 253901
rect 179969 253892 179981 253895
rect 179748 253864 179981 253892
rect 179748 253852 179754 253864
rect 179969 253861 179981 253864
rect 180015 253861 180027 253895
rect 179969 253855 180027 253861
rect 179601 253759 179659 253765
rect 179601 253725 179613 253759
rect 179647 253756 179659 253759
rect 179690 253756 179696 253768
rect 179647 253728 179696 253756
rect 179647 253725 179659 253728
rect 179601 253719 179659 253725
rect 179690 253716 179696 253728
rect 179748 253716 179754 253768
rect 336918 253172 336924 253224
rect 336976 253212 336982 253224
rect 337102 253212 337108 253224
rect 336976 253184 337108 253212
rect 336976 253172 336982 253184
rect 337102 253172 337108 253184
rect 337160 253172 337166 253224
rect 459554 253172 459560 253224
rect 459612 253212 459618 253224
rect 460474 253212 460480 253224
rect 459612 253184 460480 253212
rect 459612 253172 459618 253184
rect 460474 253172 460480 253184
rect 460532 253172 460538 253224
rect 179509 244375 179567 244381
rect 179509 244341 179521 244375
rect 179555 244372 179567 244375
rect 179690 244372 179696 244384
rect 179555 244344 179696 244372
rect 179555 244341 179567 244344
rect 179509 244335 179567 244341
rect 179690 244332 179696 244344
rect 179748 244332 179754 244384
rect 177390 244264 177396 244316
rect 177448 244304 177454 244316
rect 177448 244276 179736 244304
rect 177448 244264 177454 244276
rect 179708 244236 179736 244276
rect 177776 244208 179736 244236
rect 177776 244180 177804 244208
rect 177758 244128 177764 244180
rect 177816 244128 177822 244180
rect 179690 244128 179696 244180
rect 179748 244168 179754 244180
rect 179969 244171 180027 244177
rect 179969 244168 179981 244171
rect 179748 244140 179981 244168
rect 179748 244128 179754 244140
rect 179969 244137 179981 244140
rect 180015 244137 180027 244171
rect 179969 244131 180027 244137
rect 179598 243992 179604 244044
rect 179656 244032 179662 244044
rect 179785 244035 179843 244041
rect 179785 244032 179797 244035
rect 179656 244004 179797 244032
rect 179656 243992 179662 244004
rect 179785 244001 179797 244004
rect 179831 244001 179843 244035
rect 179785 243995 179843 244001
rect 19426 238864 19432 238876
rect 19387 238836 19432 238864
rect 19426 238824 19432 238836
rect 19484 238824 19490 238876
rect 19426 238728 19432 238740
rect 19387 238700 19432 238728
rect 19426 238688 19432 238700
rect 19484 238688 19490 238740
rect 179509 234719 179567 234725
rect 179509 234685 179521 234719
rect 179555 234716 179567 234719
rect 179598 234716 179604 234728
rect 179555 234688 179604 234716
rect 179555 234685 179567 234688
rect 179509 234679 179567 234685
rect 179598 234676 179604 234688
rect 179656 234676 179662 234728
rect 179690 234676 179696 234728
rect 179748 234716 179754 234728
rect 179969 234719 180027 234725
rect 179969 234716 179981 234719
rect 179748 234688 179981 234716
rect 179748 234676 179754 234688
rect 179969 234685 179981 234688
rect 180015 234685 180027 234719
rect 179969 234679 180027 234685
rect 179785 234651 179843 234657
rect 179785 234648 179797 234651
rect 179708 234626 179797 234648
rect 179690 234574 179696 234626
rect 179748 234620 179797 234626
rect 179748 234574 179754 234620
rect 179785 234617 179797 234620
rect 179831 234617 179843 234651
rect 179785 234611 179843 234617
rect 482094 233180 482100 233232
rect 482152 233220 482158 233232
rect 579982 233220 579988 233232
rect 482152 233192 579988 233220
rect 482152 233180 482158 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 179417 225063 179475 225069
rect 179417 225029 179429 225063
rect 179463 225060 179475 225063
rect 179598 225060 179604 225072
rect 179463 225032 179604 225060
rect 179463 225029 179475 225032
rect 179417 225023 179475 225029
rect 179598 225020 179604 225032
rect 179656 225020 179662 225072
rect 179969 224995 180027 225001
rect 179969 224992 179981 224995
rect 179616 224964 179981 224992
rect 179616 224924 179644 224964
rect 179969 224961 179981 224964
rect 180015 224961 180027 224995
rect 179969 224955 180027 224961
rect 179616 224896 179828 224924
rect 179417 224859 179475 224865
rect 179417 224825 179429 224859
rect 179463 224856 179475 224859
rect 179598 224856 179604 224868
rect 179463 224828 179604 224856
rect 179463 224825 179475 224828
rect 179417 224819 179475 224825
rect 179598 224816 179604 224828
rect 179656 224816 179662 224868
rect 179800 224856 179828 224896
rect 179969 224859 180027 224865
rect 179969 224856 179981 224859
rect 179800 224828 179981 224856
rect 179969 224825 179981 224828
rect 180015 224825 180027 224859
rect 179969 224819 180027 224825
rect 319898 223524 319904 223576
rect 319956 223564 319962 223576
rect 336918 223564 336924 223576
rect 319956 223536 336924 223564
rect 319956 223524 319962 223536
rect 336918 223524 336924 223536
rect 336976 223524 336982 223576
rect 158806 220328 158812 220380
rect 158864 220368 158870 220380
rect 160738 220368 160744 220380
rect 158864 220340 160744 220368
rect 158864 220328 158870 220340
rect 160738 220328 160744 220340
rect 160796 220328 160802 220380
rect 19426 219552 19432 219564
rect 19387 219524 19432 219552
rect 19426 219512 19432 219524
rect 19484 219512 19490 219564
rect 19426 219416 19432 219428
rect 19387 219388 19432 219416
rect 19426 219376 19432 219388
rect 19484 219376 19490 219428
rect 482186 219376 482192 219428
rect 482244 219416 482250 219428
rect 580166 219416 580172 219428
rect 482244 219388 580172 219416
rect 482244 219376 482250 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 158990 218016 158996 218068
rect 159048 218056 159054 218068
rect 160830 218056 160836 218068
rect 159048 218028 160836 218056
rect 159048 218016 159054 218028
rect 160830 218016 160836 218028
rect 160888 218016 160894 218068
rect 179414 215296 179420 215348
rect 179472 215296 179478 215348
rect 179432 215268 179460 215296
rect 179601 215271 179659 215277
rect 179601 215268 179613 215271
rect 179432 215240 179613 215268
rect 179601 215237 179613 215240
rect 179647 215237 179659 215271
rect 179601 215231 179659 215237
rect 179414 215160 179420 215212
rect 179472 215200 179478 215212
rect 179969 215203 180027 215209
rect 179969 215200 179981 215203
rect 179472 215172 179981 215200
rect 179472 215160 179478 215172
rect 179969 215169 179981 215172
rect 180015 215169 180027 215203
rect 179969 215163 180027 215169
rect 157978 211760 157984 211812
rect 158036 211800 158042 211812
rect 177022 211800 177028 211812
rect 158036 211772 177028 211800
rect 158036 211760 158042 211772
rect 177022 211760 177028 211772
rect 177080 211760 177086 211812
rect 179414 210672 179420 210724
rect 179472 210712 179478 210724
rect 179472 210684 179736 210712
rect 179472 210672 179478 210684
rect 178310 210536 178316 210588
rect 178368 210536 178374 210588
rect 179230 210536 179236 210588
rect 179288 210576 179294 210588
rect 179288 210548 179368 210576
rect 179288 210536 179294 210548
rect 178328 210372 178356 210536
rect 179340 210384 179368 210548
rect 179414 210536 179420 210588
rect 179472 210576 179478 210588
rect 179598 210576 179604 210588
rect 179472 210548 179604 210576
rect 179472 210536 179478 210548
rect 179598 210536 179604 210548
rect 179656 210536 179662 210588
rect 179708 210384 179736 210684
rect 178402 210372 178408 210384
rect 178328 210344 178408 210372
rect 178402 210332 178408 210344
rect 178460 210332 178466 210384
rect 179322 210332 179328 210384
rect 179380 210332 179386 210384
rect 179690 210332 179696 210384
rect 179748 210332 179754 210384
rect 19518 209856 19524 209908
rect 19576 209896 19582 209908
rect 19613 209899 19671 209905
rect 19613 209896 19625 209899
rect 19576 209868 19625 209896
rect 19576 209856 19582 209868
rect 19613 209865 19625 209868
rect 19659 209865 19671 209899
rect 19613 209859 19671 209865
rect 19981 209831 20039 209837
rect 19981 209828 19993 209831
rect 19628 209800 19993 209828
rect 19426 209760 19432 209772
rect 19387 209732 19432 209760
rect 19426 209720 19432 209732
rect 19484 209720 19490 209772
rect 19628 209760 19656 209800
rect 19981 209797 19993 209800
rect 20027 209797 20039 209831
rect 19981 209791 20039 209797
rect 19628 209732 19748 209760
rect 19518 209692 19524 209704
rect 19479 209664 19524 209692
rect 19518 209652 19524 209664
rect 19576 209652 19582 209704
rect 19518 209516 19524 209568
rect 19576 209556 19582 209568
rect 19720 209556 19748 209732
rect 19794 209720 19800 209772
rect 19852 209720 19858 209772
rect 19576 209528 19748 209556
rect 19576 209516 19582 209528
rect 19426 209448 19432 209500
rect 19484 209488 19490 209500
rect 19812 209488 19840 209720
rect 19484 209460 19840 209488
rect 19484 209448 19490 209460
rect 19610 209420 19616 209432
rect 19571 209392 19616 209420
rect 19610 209380 19616 209392
rect 19668 209380 19674 209432
rect 19521 209355 19579 209361
rect 19521 209321 19533 209355
rect 19567 209352 19579 209355
rect 19794 209352 19800 209364
rect 19567 209324 19800 209352
rect 19567 209321 19579 209324
rect 19521 209315 19579 209321
rect 19794 209312 19800 209324
rect 19852 209312 19858 209364
rect 178402 205912 178408 205964
rect 178460 205912 178466 205964
rect 178494 205912 178500 205964
rect 178552 205912 178558 205964
rect 178586 205912 178592 205964
rect 178644 205912 178650 205964
rect 179322 205952 179328 205964
rect 178696 205924 179328 205952
rect 178034 205748 178040 205760
rect 177995 205720 178040 205748
rect 178034 205708 178040 205720
rect 178092 205708 178098 205760
rect 178420 205680 178448 205912
rect 178512 205692 178540 205912
rect 178604 205692 178632 205912
rect 178696 205692 178724 205924
rect 179322 205912 179328 205924
rect 179380 205912 179386 205964
rect 179690 205816 179696 205828
rect 179651 205788 179696 205816
rect 179690 205776 179696 205788
rect 179748 205776 179754 205828
rect 178144 205652 178448 205680
rect 178034 205572 178040 205624
rect 178092 205612 178098 205624
rect 178144 205612 178172 205652
rect 178494 205640 178500 205692
rect 178552 205640 178558 205692
rect 178586 205640 178592 205692
rect 178644 205640 178650 205692
rect 178678 205640 178684 205692
rect 178736 205640 178742 205692
rect 179601 205683 179659 205689
rect 179601 205649 179613 205683
rect 179647 205680 179659 205683
rect 179690 205680 179696 205692
rect 179647 205652 179696 205680
rect 179647 205649 179659 205652
rect 179601 205643 179659 205649
rect 179690 205640 179696 205652
rect 179748 205640 179754 205692
rect 178092 205584 178172 205612
rect 178092 205572 178098 205584
rect 165801 204323 165859 204329
rect 165801 204289 165813 204323
rect 165847 204320 165859 204323
rect 165847 204292 166580 204320
rect 165847 204289 165859 204292
rect 165801 204283 165859 204289
rect 159358 204212 159364 204264
rect 159416 204252 159422 204264
rect 165985 204255 166043 204261
rect 165985 204252 165997 204255
rect 159416 204224 165997 204252
rect 159416 204212 159422 204224
rect 165985 204221 165997 204224
rect 166031 204221 166043 204255
rect 165985 204215 166043 204221
rect 166077 204255 166135 204261
rect 166077 204221 166089 204255
rect 166123 204252 166135 204255
rect 166552 204252 166580 204292
rect 177482 204252 177488 204264
rect 166123 204224 166488 204252
rect 166552 204224 177488 204252
rect 166123 204221 166135 204224
rect 166077 204215 166135 204221
rect 160738 204144 160744 204196
rect 160796 204184 160802 204196
rect 165893 204187 165951 204193
rect 165893 204184 165905 204187
rect 160796 204156 165905 204184
rect 160796 204144 160802 204156
rect 165893 204153 165905 204156
rect 165939 204153 165951 204187
rect 165893 204147 165951 204153
rect 166169 204187 166227 204193
rect 166169 204153 166181 204187
rect 166215 204184 166227 204187
rect 166460 204184 166488 204224
rect 177482 204212 177488 204224
rect 177540 204212 177546 204264
rect 177574 204184 177580 204196
rect 166215 204156 166396 204184
rect 166460 204156 177580 204184
rect 166215 204153 166227 204156
rect 166169 204147 166227 204153
rect 160830 204076 160836 204128
rect 160888 204116 160894 204128
rect 166368 204116 166396 204156
rect 177574 204144 177580 204156
rect 177632 204144 177638 204196
rect 175737 204119 175795 204125
rect 175737 204116 175749 204119
rect 160888 204088 166304 204116
rect 166368 204088 175749 204116
rect 160888 204076 160894 204088
rect 17494 204008 17500 204060
rect 17552 204048 17558 204060
rect 166169 204051 166227 204057
rect 166169 204048 166181 204051
rect 17552 204020 166181 204048
rect 17552 204008 17558 204020
rect 166169 204017 166181 204020
rect 166215 204017 166227 204051
rect 166276 204048 166304 204088
rect 175737 204085 175749 204088
rect 175783 204085 175795 204119
rect 175737 204079 175795 204085
rect 176105 204119 176163 204125
rect 176105 204085 176117 204119
rect 176151 204116 176163 204119
rect 177666 204116 177672 204128
rect 176151 204088 177672 204116
rect 176151 204085 176163 204088
rect 176105 204079 176163 204085
rect 177666 204076 177672 204088
rect 177724 204076 177730 204128
rect 175921 204051 175979 204057
rect 166276 204020 175780 204048
rect 166169 204011 166227 204017
rect 17402 203940 17408 203992
rect 17460 203980 17466 203992
rect 166077 203983 166135 203989
rect 166077 203980 166089 203983
rect 17460 203952 166089 203980
rect 17460 203940 17466 203952
rect 166077 203949 166089 203952
rect 166123 203949 166135 203983
rect 175645 203983 175703 203989
rect 175645 203980 175657 203983
rect 166077 203943 166135 203949
rect 166276 203952 175657 203980
rect 19429 203915 19487 203921
rect 19429 203881 19441 203915
rect 19475 203912 19487 203915
rect 20070 203912 20076 203924
rect 19475 203884 20076 203912
rect 19475 203881 19487 203884
rect 19429 203875 19487 203881
rect 20070 203872 20076 203884
rect 20128 203872 20134 203924
rect 159542 203872 159548 203924
rect 159600 203912 159606 203924
rect 166276 203912 166304 203952
rect 175645 203949 175657 203952
rect 175691 203949 175703 203983
rect 175752 203980 175780 204020
rect 175921 204017 175933 204051
rect 175967 204048 175979 204051
rect 181625 204051 181683 204057
rect 175967 204020 181576 204048
rect 175967 204017 175979 204020
rect 175921 204011 175979 204017
rect 181441 203983 181499 203989
rect 181441 203980 181453 203983
rect 175752 203952 181453 203980
rect 175645 203943 175703 203949
rect 181441 203949 181453 203952
rect 181487 203949 181499 203983
rect 181548 203980 181576 204020
rect 181625 204017 181637 204051
rect 181671 204048 181683 204051
rect 318886 204048 318892 204060
rect 181671 204020 318892 204048
rect 181671 204017 181683 204020
rect 181625 204011 181683 204017
rect 318886 204008 318892 204020
rect 318944 204008 318950 204060
rect 317598 203980 317604 203992
rect 181548 203952 317604 203980
rect 181441 203943 181499 203949
rect 317598 203940 317604 203952
rect 317656 203940 317662 203992
rect 317414 203912 317420 203924
rect 159600 203884 166304 203912
rect 166368 203884 317420 203912
rect 159600 203872 159606 203884
rect 17678 203804 17684 203856
rect 17736 203844 17742 203856
rect 165801 203847 165859 203853
rect 165801 203844 165813 203847
rect 17736 203816 165813 203844
rect 17736 203804 17742 203816
rect 165801 203813 165813 203816
rect 165847 203813 165859 203847
rect 165801 203807 165859 203813
rect 165985 203847 166043 203853
rect 165985 203813 165997 203847
rect 166031 203844 166043 203847
rect 166368 203844 166396 203884
rect 317414 203872 317420 203884
rect 317472 203872 317478 203924
rect 166031 203816 166396 203844
rect 166445 203847 166503 203853
rect 166031 203813 166043 203816
rect 165985 203807 166043 203813
rect 166445 203813 166457 203847
rect 166491 203844 166503 203847
rect 318794 203844 318800 203856
rect 166491 203816 318800 203844
rect 166491 203813 166503 203816
rect 166445 203807 166503 203813
rect 318794 203804 318800 203816
rect 318852 203804 318858 203856
rect 3602 203736 3608 203788
rect 3660 203776 3666 203788
rect 331950 203776 331956 203788
rect 3660 203748 331956 203776
rect 3660 203736 3666 203748
rect 331950 203736 331956 203748
rect 332008 203736 332014 203788
rect 30282 203668 30288 203720
rect 30340 203708 30346 203720
rect 370498 203708 370504 203720
rect 30340 203680 370504 203708
rect 30340 203668 30346 203680
rect 370498 203668 370504 203680
rect 370556 203668 370562 203720
rect 27522 203600 27528 203652
rect 27580 203640 27586 203652
rect 367738 203640 367744 203652
rect 27580 203612 367744 203640
rect 27580 203600 27586 203612
rect 367738 203600 367744 203612
rect 367796 203600 367802 203652
rect 106182 203532 106188 203584
rect 106240 203572 106246 203584
rect 458174 203572 458180 203584
rect 106240 203544 458180 203572
rect 106240 203532 106246 203544
rect 458174 203532 458180 203544
rect 458232 203532 458238 203584
rect 17770 203464 17776 203516
rect 17828 203504 17834 203516
rect 166169 203507 166227 203513
rect 166169 203504 166181 203507
rect 17828 203476 166181 203504
rect 17828 203464 17834 203476
rect 166169 203473 166181 203476
rect 166215 203473 166227 203507
rect 166169 203467 166227 203473
rect 166261 203507 166319 203513
rect 166261 203473 166273 203507
rect 166307 203504 166319 203507
rect 317506 203504 317512 203516
rect 166307 203476 317512 203504
rect 166307 203473 166319 203476
rect 166261 203467 166319 203473
rect 317506 203464 317512 203476
rect 317564 203464 317570 203516
rect 17586 203396 17592 203448
rect 17644 203436 17650 203448
rect 177758 203436 177764 203448
rect 17644 203408 177764 203436
rect 17644 203396 17650 203408
rect 177758 203396 177764 203408
rect 177816 203396 177822 203448
rect 179506 203396 179512 203448
rect 179564 203436 179570 203448
rect 179564 203408 186314 203436
rect 179564 203396 179570 203408
rect 16666 203328 16672 203380
rect 16724 203368 16730 203380
rect 69750 203368 69756 203380
rect 16724 203340 69756 203368
rect 16724 203328 16730 203340
rect 69750 203328 69756 203340
rect 69808 203328 69814 203380
rect 159450 203328 159456 203380
rect 159508 203368 159514 203380
rect 166261 203371 166319 203377
rect 166261 203368 166273 203371
rect 159508 203340 166273 203368
rect 159508 203328 159514 203340
rect 166261 203337 166273 203340
rect 166307 203337 166319 203371
rect 166261 203331 166319 203337
rect 176470 203328 176476 203380
rect 176528 203368 176534 203380
rect 186286 203368 186314 203408
rect 231118 203368 231124 203380
rect 176528 203340 181484 203368
rect 186286 203340 231124 203368
rect 176528 203328 176534 203340
rect 17310 203260 17316 203312
rect 17368 203300 17374 203312
rect 71130 203300 71136 203312
rect 17368 203272 71136 203300
rect 17368 203260 17374 203272
rect 71130 203260 71136 203272
rect 71188 203260 71194 203312
rect 166169 203303 166227 203309
rect 166169 203269 166181 203303
rect 166215 203300 166227 203303
rect 177390 203300 177396 203312
rect 166215 203272 177396 203300
rect 166215 203269 166227 203272
rect 166169 203263 166227 203269
rect 177390 203260 177396 203272
rect 177448 203260 177454 203312
rect 179693 203303 179751 203309
rect 179693 203269 179705 203303
rect 179739 203300 179751 203303
rect 180058 203300 180064 203312
rect 179739 203272 180064 203300
rect 179739 203269 179751 203272
rect 179693 203263 179751 203269
rect 180058 203260 180064 203272
rect 180116 203260 180122 203312
rect 181456 203300 181484 203340
rect 231118 203328 231124 203340
rect 231176 203328 231182 203380
rect 229738 203300 229744 203312
rect 181456 203272 229744 203300
rect 229738 203260 229744 203272
rect 229796 203260 229802 203312
rect 18230 203192 18236 203244
rect 18288 203232 18294 203244
rect 72234 203232 72240 203244
rect 18288 203204 72240 203232
rect 18288 203192 18294 203204
rect 72234 203192 72240 203204
rect 72292 203192 72298 203244
rect 178494 203192 178500 203244
rect 178552 203232 178558 203244
rect 232222 203232 232228 203244
rect 178552 203204 232228 203232
rect 178552 203192 178558 203204
rect 232222 203192 232228 203204
rect 232280 203192 232286 203244
rect 19610 203124 19616 203176
rect 19668 203164 19674 203176
rect 75730 203164 75736 203176
rect 19668 203136 75736 203164
rect 19668 203124 19674 203136
rect 75730 203124 75736 203136
rect 75788 203124 75794 203176
rect 179598 203124 179604 203176
rect 179656 203164 179662 203176
rect 233326 203164 233332 203176
rect 179656 203136 233332 203164
rect 179656 203124 179662 203136
rect 233326 203124 233332 203136
rect 233384 203124 233390 203176
rect 18138 203056 18144 203108
rect 18196 203096 18202 203108
rect 73338 203096 73344 203108
rect 18196 203068 73344 203096
rect 18196 203056 18202 203068
rect 73338 203056 73344 203068
rect 73396 203056 73402 203108
rect 178037 203099 178095 203105
rect 178037 203065 178049 203099
rect 178083 203096 178095 203099
rect 178494 203096 178500 203108
rect 178083 203068 178500 203096
rect 178083 203065 178095 203068
rect 178037 203059 178095 203065
rect 178494 203056 178500 203068
rect 178552 203056 178558 203108
rect 179414 203056 179420 203108
rect 179472 203096 179478 203108
rect 234430 203096 234436 203108
rect 179472 203068 234436 203096
rect 179472 203056 179478 203068
rect 234430 203056 234436 203068
rect 234488 203056 234494 203108
rect 17954 202988 17960 203040
rect 18012 203028 18018 203040
rect 74350 203028 74356 203040
rect 18012 203000 74356 203028
rect 18012 202988 18018 203000
rect 74350 202988 74356 203000
rect 74408 202988 74414 203040
rect 179690 202988 179696 203040
rect 179748 203028 179754 203040
rect 235718 203028 235724 203040
rect 179748 203000 235724 203028
rect 179748 202988 179754 203000
rect 235718 202988 235724 203000
rect 235776 202988 235782 203040
rect 17218 202920 17224 202972
rect 17276 202960 17282 202972
rect 76926 202960 76932 202972
rect 17276 202932 76932 202960
rect 17276 202920 17282 202932
rect 76926 202920 76932 202932
rect 76984 202920 76990 202972
rect 177942 202920 177948 202972
rect 178000 202960 178006 202972
rect 238018 202960 238024 202972
rect 178000 202932 238024 202960
rect 178000 202920 178006 202932
rect 238018 202920 238024 202932
rect 238076 202920 238082 202972
rect 17126 202852 17132 202904
rect 17184 202892 17190 202904
rect 78030 202892 78036 202904
rect 17184 202864 78036 202892
rect 17184 202852 17190 202864
rect 78030 202852 78036 202864
rect 78088 202852 78094 202904
rect 176378 202852 176384 202904
rect 176436 202892 176442 202904
rect 237006 202892 237012 202904
rect 176436 202864 237012 202892
rect 176436 202852 176442 202864
rect 237006 202852 237012 202864
rect 237064 202852 237070 202904
rect 17862 202784 17868 202836
rect 17920 202824 17926 202836
rect 157978 202824 157984 202836
rect 17920 202796 157984 202824
rect 17920 202784 17926 202796
rect 157978 202784 157984 202796
rect 158036 202784 158042 202836
rect 3510 202716 3516 202768
rect 3568 202756 3574 202768
rect 334710 202756 334716 202768
rect 3568 202728 334716 202756
rect 3568 202716 3574 202728
rect 334710 202716 334716 202728
rect 334768 202716 334774 202768
rect 119890 202240 119896 202292
rect 119948 202280 119954 202292
rect 436738 202280 436744 202292
rect 119948 202252 436744 202280
rect 119948 202240 119954 202252
rect 436738 202240 436744 202252
rect 436796 202240 436802 202292
rect 23382 202172 23388 202224
rect 23440 202212 23446 202224
rect 347038 202212 347044 202224
rect 23440 202184 347044 202212
rect 23440 202172 23446 202184
rect 347038 202172 347044 202184
rect 347096 202172 347102 202224
rect 113082 202104 113088 202156
rect 113140 202144 113146 202156
rect 465074 202144 465080 202156
rect 113140 202116 465080 202144
rect 113140 202104 113146 202116
rect 465074 202104 465080 202116
rect 465132 202104 465138 202156
rect 17218 201968 17224 202020
rect 17276 202008 17282 202020
rect 17862 202008 17868 202020
rect 17276 201980 17868 202008
rect 17276 201968 17282 201980
rect 17862 201968 17868 201980
rect 17920 201968 17926 202020
rect 19702 201424 19708 201476
rect 19760 201464 19766 201476
rect 67634 201464 67640 201476
rect 19760 201436 67640 201464
rect 19760 201424 19766 201436
rect 67634 201424 67640 201436
rect 67692 201424 67698 201476
rect 79962 201424 79968 201476
rect 80020 201464 80026 201476
rect 157334 201464 157340 201476
rect 80020 201436 157340 201464
rect 80020 201424 80026 201436
rect 157334 201424 157340 201436
rect 157392 201424 157398 201476
rect 179782 201424 179788 201476
rect 179840 201464 179846 201476
rect 224954 201464 224960 201476
rect 179840 201436 224960 201464
rect 179840 201424 179846 201436
rect 224954 201424 224960 201436
rect 225012 201424 225018 201476
rect 238938 201424 238944 201476
rect 238996 201464 239002 201476
rect 316586 201464 316592 201476
rect 238996 201436 316592 201464
rect 238996 201424 239002 201436
rect 316586 201424 316592 201436
rect 316644 201424 316650 201476
rect 19518 201356 19524 201408
rect 19576 201396 19582 201408
rect 37274 201396 37280 201408
rect 19576 201368 37280 201396
rect 19576 201356 19582 201368
rect 37274 201356 37280 201368
rect 37332 201356 37338 201408
rect 179874 201356 179880 201408
rect 179932 201396 179938 201408
rect 223574 201396 223580 201408
rect 179932 201368 223580 201396
rect 179932 201356 179938 201368
rect 223574 201356 223580 201368
rect 223632 201356 223638 201408
rect 302234 201356 302240 201408
rect 302292 201396 302298 201408
rect 303154 201396 303160 201408
rect 302292 201368 303160 201396
rect 302292 201356 302298 201368
rect 303154 201356 303160 201368
rect 303212 201396 303218 201408
rect 336826 201396 336832 201408
rect 303212 201368 336832 201396
rect 303212 201356 303218 201368
rect 336826 201356 336832 201368
rect 336884 201356 336890 201408
rect 19334 201288 19340 201340
rect 19392 201328 19398 201340
rect 36538 201328 36544 201340
rect 19392 201300 36544 201328
rect 19392 201288 19398 201300
rect 36538 201288 36544 201300
rect 36596 201288 36602 201340
rect 179966 201288 179972 201340
rect 180024 201328 180030 201340
rect 222194 201328 222200 201340
rect 180024 201300 222200 201328
rect 180024 201288 180030 201300
rect 222194 201288 222200 201300
rect 222252 201288 222258 201340
rect 302326 201288 302332 201340
rect 302384 201328 302390 201340
rect 303522 201328 303528 201340
rect 302384 201300 303528 201328
rect 302384 201288 302390 201300
rect 303522 201288 303528 201300
rect 303580 201328 303586 201340
rect 337010 201328 337016 201340
rect 303580 201300 337016 201328
rect 303580 201288 303586 201300
rect 337010 201288 337016 201300
rect 337068 201288 337074 201340
rect 19978 201220 19984 201272
rect 20036 201260 20042 201272
rect 63494 201260 63500 201272
rect 20036 201232 63500 201260
rect 20036 201220 20042 201232
rect 63494 201220 63500 201232
rect 63552 201220 63558 201272
rect 180058 201220 180064 201272
rect 180116 201260 180122 201272
rect 195974 201260 195980 201272
rect 180116 201232 195980 201260
rect 180116 201220 180122 201232
rect 195974 201220 195980 201232
rect 196032 201220 196038 201272
rect 19242 201152 19248 201204
rect 19300 201192 19306 201204
rect 62114 201192 62120 201204
rect 19300 201164 62120 201192
rect 19300 201152 19306 201164
rect 62114 201152 62120 201164
rect 62172 201152 62178 201204
rect 179138 201152 179144 201204
rect 179196 201192 179202 201204
rect 219986 201192 219992 201204
rect 179196 201164 219992 201192
rect 179196 201152 179202 201164
rect 219986 201152 219992 201164
rect 220044 201152 220050 201204
rect 18414 201084 18420 201136
rect 18472 201124 18478 201136
rect 59354 201124 59360 201136
rect 18472 201096 59360 201124
rect 18472 201084 18478 201096
rect 59354 201084 59360 201096
rect 59412 201084 59418 201136
rect 179230 201084 179236 201136
rect 179288 201124 179294 201136
rect 219434 201124 219440 201136
rect 179288 201096 219440 201124
rect 179288 201084 179294 201096
rect 219434 201084 219440 201096
rect 219492 201084 219498 201136
rect 18966 201016 18972 201068
rect 19024 201056 19030 201068
rect 59446 201056 59452 201068
rect 19024 201028 59452 201056
rect 19024 201016 19030 201028
rect 59446 201016 59452 201028
rect 59504 201016 59510 201068
rect 179046 201016 179052 201068
rect 179104 201056 179110 201068
rect 215294 201056 215300 201068
rect 179104 201028 215300 201056
rect 179104 201016 179110 201028
rect 215294 201016 215300 201028
rect 215352 201016 215358 201068
rect 18690 200948 18696 201000
rect 18748 200988 18754 201000
rect 55582 200988 55588 201000
rect 18748 200960 55588 200988
rect 18748 200948 18754 200960
rect 55582 200948 55588 200960
rect 55640 200948 55646 201000
rect 178586 200948 178592 201000
rect 178644 200988 178650 201000
rect 211154 200988 211160 201000
rect 178644 200960 211160 200988
rect 178644 200948 178650 200960
rect 211154 200948 211160 200960
rect 211212 200948 211218 201000
rect 19794 200880 19800 200932
rect 19852 200920 19858 200932
rect 52454 200920 52460 200932
rect 19852 200892 52460 200920
rect 19852 200880 19858 200892
rect 52454 200880 52460 200892
rect 52512 200880 52518 200932
rect 143442 200880 143448 200932
rect 143500 200920 143506 200932
rect 302234 200920 302240 200932
rect 143500 200892 302240 200920
rect 143500 200880 143506 200892
rect 302234 200880 302240 200892
rect 302292 200880 302298 200932
rect 18506 200812 18512 200864
rect 18564 200852 18570 200864
rect 51074 200852 51080 200864
rect 18564 200824 51080 200852
rect 18564 200812 18570 200824
rect 51074 200812 51080 200824
rect 51132 200812 51138 200864
rect 178862 200812 178868 200864
rect 178920 200852 178926 200864
rect 211246 200852 211252 200864
rect 178920 200824 211252 200852
rect 178920 200812 178926 200824
rect 211246 200812 211252 200824
rect 211304 200812 211310 200864
rect 18598 200744 18604 200796
rect 18656 200784 18662 200796
rect 51166 200784 51172 200796
rect 18656 200756 51172 200784
rect 18656 200744 18662 200756
rect 51166 200744 51172 200756
rect 51224 200744 51230 200796
rect 143442 200744 143448 200796
rect 143500 200784 143506 200796
rect 302326 200784 302332 200796
rect 143500 200756 302332 200784
rect 143500 200744 143506 200756
rect 302326 200744 302332 200756
rect 302384 200744 302390 200796
rect 19058 200676 19064 200728
rect 19116 200716 19122 200728
rect 49694 200716 49700 200728
rect 19116 200688 49700 200716
rect 19116 200676 19122 200688
rect 49694 200676 49700 200688
rect 49752 200676 49758 200728
rect 178770 200676 178776 200728
rect 178828 200716 178834 200728
rect 209866 200716 209872 200728
rect 178828 200688 209872 200716
rect 178828 200676 178834 200688
rect 209866 200676 209872 200688
rect 209924 200676 209930 200728
rect 18322 200608 18328 200660
rect 18380 200648 18386 200660
rect 44358 200648 44364 200660
rect 18380 200620 44364 200648
rect 18380 200608 18386 200620
rect 44358 200608 44364 200620
rect 44416 200608 44422 200660
rect 178126 200608 178132 200660
rect 178184 200648 178190 200660
rect 204346 200648 204352 200660
rect 178184 200620 204352 200648
rect 178184 200608 178190 200620
rect 204346 200608 204352 200620
rect 204404 200608 204410 200660
rect 18874 200540 18880 200592
rect 18932 200580 18938 200592
rect 44174 200580 44180 200592
rect 18932 200552 44180 200580
rect 18932 200540 18938 200552
rect 44174 200540 44180 200552
rect 44232 200540 44238 200592
rect 178218 200540 178224 200592
rect 178276 200580 178282 200592
rect 204254 200580 204260 200592
rect 178276 200552 204260 200580
rect 178276 200540 178282 200552
rect 204254 200540 204260 200552
rect 204312 200540 204318 200592
rect 18046 200472 18052 200524
rect 18104 200512 18110 200524
rect 41598 200512 41604 200524
rect 18104 200484 41604 200512
rect 18104 200472 18110 200484
rect 41598 200472 41604 200484
rect 41656 200472 41662 200524
rect 176562 200472 176568 200524
rect 176620 200512 176626 200524
rect 200114 200512 200120 200524
rect 176620 200484 200120 200512
rect 176620 200472 176626 200484
rect 200114 200472 200120 200484
rect 200172 200472 200178 200524
rect 20070 200404 20076 200456
rect 20128 200444 20134 200456
rect 40034 200444 40040 200456
rect 20128 200416 40040 200444
rect 20128 200404 20134 200416
rect 40034 200404 40040 200416
rect 40092 200404 40098 200456
rect 178402 200404 178408 200456
rect 178460 200444 178466 200456
rect 201494 200444 201500 200456
rect 178460 200416 201500 200444
rect 178460 200404 178466 200416
rect 201494 200404 201500 200416
rect 201552 200404 201558 200456
rect 18782 200336 18788 200388
rect 18840 200376 18846 200388
rect 38654 200376 38660 200388
rect 18840 200348 38660 200376
rect 18840 200336 18846 200348
rect 38654 200336 38660 200348
rect 38712 200336 38718 200388
rect 178310 200336 178316 200388
rect 178368 200376 178374 200388
rect 198734 200376 198740 200388
rect 178368 200348 198740 200376
rect 178368 200336 178374 200348
rect 198734 200336 198740 200348
rect 198792 200336 198798 200388
rect 19886 200268 19892 200320
rect 19944 200308 19950 200320
rect 66254 200308 66260 200320
rect 19944 200280 66260 200308
rect 19944 200268 19950 200280
rect 66254 200268 66260 200280
rect 66312 200268 66318 200320
rect 178034 200268 178040 200320
rect 178092 200308 178098 200320
rect 197354 200308 197360 200320
rect 178092 200280 197360 200308
rect 178092 200268 178098 200280
rect 197354 200268 197360 200280
rect 197412 200268 197418 200320
rect 19150 200200 19156 200252
rect 19208 200240 19214 200252
rect 64874 200240 64880 200252
rect 19208 200212 64880 200240
rect 19208 200200 19214 200212
rect 64874 200200 64880 200212
rect 64932 200200 64938 200252
rect 178494 200200 178500 200252
rect 178552 200240 178558 200252
rect 196158 200240 196164 200252
rect 178552 200212 196164 200240
rect 178552 200200 178558 200212
rect 196158 200200 196164 200212
rect 196216 200200 196222 200252
rect 201126 200200 201132 200252
rect 201184 200240 201190 200252
rect 201862 200240 201868 200252
rect 201184 200212 201868 200240
rect 201184 200200 201190 200212
rect 201862 200200 201868 200212
rect 201920 200200 201926 200252
rect 19426 200132 19432 200184
rect 19484 200172 19490 200184
rect 35894 200172 35900 200184
rect 19484 200144 35900 200172
rect 19484 200132 19490 200144
rect 35894 200132 35900 200144
rect 35952 200132 35958 200184
rect 178678 200132 178684 200184
rect 178736 200172 178742 200184
rect 220814 200172 220820 200184
rect 178736 200144 220820 200172
rect 178736 200132 178742 200144
rect 220814 200132 220820 200144
rect 220872 200132 220878 200184
rect 482922 193128 482928 193180
rect 482980 193168 482986 193180
rect 580166 193168 580172 193180
rect 482980 193140 580172 193168
rect 482980 193128 482986 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3602 188300 3608 188352
rect 3660 188340 3666 188352
rect 330478 188340 330484 188352
rect 3660 188312 330484 188340
rect 3660 188300 3666 188312
rect 330478 188300 330484 188312
rect 330536 188300 330542 188352
rect 482830 179324 482836 179376
rect 482888 179364 482894 179376
rect 580166 179364 580172 179376
rect 482888 179336 580172 179364
rect 482888 179324 482894 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 482738 153144 482744 153196
rect 482796 153184 482802 153196
rect 580166 153184 580172 153196
rect 482796 153156 580172 153184
rect 482796 153144 482802 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 325050 150396 325056 150408
rect 3384 150368 325056 150396
rect 3384 150356 3390 150368
rect 325050 150356 325056 150368
rect 325108 150356 325114 150408
rect 482646 139340 482652 139392
rect 482704 139380 482710 139392
rect 580166 139380 580172 139392
rect 482704 139352 580172 139380
rect 482704 139340 482710 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137232 3516 137284
rect 3568 137272 3574 137284
rect 329098 137272 329104 137284
rect 3568 137244 329104 137272
rect 3568 137232 3574 137244
rect 329098 137232 329104 137244
rect 329156 137232 329162 137284
rect 482554 113092 482560 113144
rect 482612 113132 482618 113144
rect 579798 113132 579804 113144
rect 482612 113104 579804 113132
rect 482612 113092 482618 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 482462 100648 482468 100700
rect 482520 100688 482526 100700
rect 580166 100688 580172 100700
rect 482520 100660 580172 100688
rect 482520 100648 482526 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 323578 97968 323584 97980
rect 3292 97940 323584 97968
rect 3292 97928 3298 97940
rect 323578 97928 323584 97940
rect 323636 97928 323642 97980
rect 3602 84804 3608 84856
rect 3660 84844 3666 84856
rect 335998 84844 336004 84856
rect 3660 84816 336004 84844
rect 3660 84804 3666 84816
rect 335998 84804 336004 84816
rect 336056 84804 336062 84856
rect 485038 73108 485044 73160
rect 485096 73148 485102 73160
rect 580166 73148 580172 73160
rect 485096 73120 580172 73148
rect 485096 73108 485102 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 482370 60664 482376 60716
rect 482428 60704 482434 60716
rect 580166 60704 580172 60716
rect 482428 60676 580172 60704
rect 482428 60664 482434 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 32398 51824 32404 51876
rect 32456 51864 32462 51876
rect 369854 51864 369860 51876
rect 32456 51836 369860 51864
rect 32456 51824 32462 51836
rect 369854 51824 369860 51836
rect 369912 51824 369918 51876
rect 43438 51756 43444 51808
rect 43496 51796 43502 51808
rect 382274 51796 382280 51808
rect 43496 51768 382280 51796
rect 43496 51756 43502 51768
rect 382274 51756 382280 51768
rect 382332 51756 382338 51808
rect 35158 51688 35164 51740
rect 35216 51728 35222 51740
rect 373994 51728 374000 51740
rect 35216 51700 374000 51728
rect 35216 51688 35222 51700
rect 373994 51688 374000 51700
rect 374052 51688 374058 51740
rect 3418 44820 3424 44872
rect 3476 44860 3482 44872
rect 320818 44860 320824 44872
rect 3476 44832 320824 44860
rect 3476 44820 3482 44832
rect 320818 44820 320824 44832
rect 320876 44820 320882 44872
rect 483658 33056 483664 33108
rect 483716 33096 483722 33108
rect 580166 33096 580172 33108
rect 483716 33068 580172 33096
rect 483716 33056 483722 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 34422 29860 34428 29912
rect 34480 29900 34486 29912
rect 376754 29900 376760 29912
rect 34480 29872 376760 29900
rect 34480 29860 34486 29872
rect 376754 29860 376760 29872
rect 376812 29860 376818 29912
rect 41322 29792 41328 29844
rect 41380 29832 41386 29844
rect 385034 29832 385040 29844
rect 41380 29804 385040 29832
rect 41380 29792 41386 29804
rect 385034 29792 385040 29804
rect 385092 29792 385098 29844
rect 37182 29724 37188 29776
rect 37240 29764 37246 29776
rect 380894 29764 380900 29776
rect 37240 29736 380900 29764
rect 37240 29724 37246 29736
rect 380894 29724 380900 29736
rect 380952 29724 380958 29776
rect 55122 29656 55128 29708
rect 55180 29696 55186 29708
rect 400214 29696 400220 29708
rect 55180 29668 400220 29696
rect 55180 29656 55186 29668
rect 400214 29656 400220 29668
rect 400272 29656 400278 29708
rect 48222 29588 48228 29640
rect 48280 29628 48286 29640
rect 393314 29628 393320 29640
rect 48280 29600 393320 29628
rect 48280 29588 48286 29600
rect 393314 29588 393320 29600
rect 393372 29588 393378 29640
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 322198 20652 322204 20664
rect 3568 20624 322204 20652
rect 3568 20612 3574 20624
rect 322198 20612 322204 20624
rect 322256 20612 322262 20664
rect 482278 20612 482284 20664
rect 482336 20652 482342 20664
rect 579982 20652 579988 20664
rect 482336 20624 579988 20652
rect 482336 20612 482342 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 59262 13268 59268 13320
rect 59320 13308 59326 13320
rect 318058 13308 318064 13320
rect 59320 13280 318064 13308
rect 59320 13268 59326 13280
rect 318058 13268 318064 13280
rect 318116 13268 318122 13320
rect 52362 13200 52368 13252
rect 52420 13240 52426 13252
rect 340230 13240 340236 13252
rect 52420 13212 340236 13240
rect 52420 13200 52426 13212
rect 340230 13200 340236 13212
rect 340288 13200 340294 13252
rect 22738 13132 22744 13184
rect 22796 13172 22802 13184
rect 360194 13172 360200 13184
rect 22796 13144 360200 13172
rect 22796 13132 22802 13144
rect 360194 13132 360200 13144
rect 360252 13132 360258 13184
rect 39298 13064 39304 13116
rect 39356 13104 39362 13116
rect 378134 13104 378140 13116
rect 39356 13076 378140 13104
rect 39356 13064 39362 13076
rect 378134 13064 378140 13076
rect 378192 13064 378198 13116
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 342254 11744 342260 11756
rect 14516 11716 342260 11744
rect 14516 11704 14522 11716
rect 342254 11704 342260 11716
rect 342312 11704 342318 11756
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 349154 10520 349160 10532
rect 18656 10492 349160 10520
rect 18656 10480 18662 10492
rect 349154 10480 349160 10492
rect 349212 10480 349218 10532
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 340874 10452 340880 10464
rect 7616 10424 340880 10452
rect 7616 10412 7622 10424
rect 340874 10412 340880 10424
rect 340932 10412 340938 10464
rect 66162 10344 66168 10396
rect 66220 10384 66226 10396
rect 412634 10384 412640 10396
rect 66220 10356 412640 10384
rect 66220 10344 66226 10356
rect 412634 10344 412640 10356
rect 412692 10344 412698 10396
rect 124122 10276 124128 10328
rect 124180 10316 124186 10328
rect 475378 10316 475384 10328
rect 124180 10288 475384 10316
rect 124180 10276 124186 10288
rect 475378 10276 475384 10288
rect 475436 10276 475442 10328
rect 9950 9188 9956 9240
rect 10008 9228 10014 9240
rect 320910 9228 320916 9240
rect 10008 9200 320916 9228
rect 10008 9188 10014 9200
rect 320910 9188 320916 9200
rect 320968 9188 320974 9240
rect 45462 9120 45468 9172
rect 45520 9160 45526 9172
rect 374638 9160 374644 9172
rect 45520 9132 374644 9160
rect 45520 9120 45526 9132
rect 374638 9120 374644 9132
rect 374696 9120 374702 9172
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 340138 9092 340144 9104
rect 4120 9064 340144 9092
rect 4120 9052 4126 9064
rect 340138 9052 340144 9064
rect 340196 9052 340202 9104
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 345658 9024 345664 9036
rect 7708 8996 345664 9024
rect 7708 8984 7714 8996
rect 345658 8984 345664 8996
rect 345716 8984 345722 9036
rect 44266 8916 44272 8968
rect 44324 8956 44330 8968
rect 389174 8956 389180 8968
rect 44324 8928 389180 8956
rect 44324 8916 44330 8928
rect 389174 8916 389180 8928
rect 389232 8916 389238 8968
rect 71498 8236 71504 8288
rect 71556 8276 71562 8288
rect 419534 8276 419540 8288
rect 71556 8248 419540 8276
rect 71556 8236 71562 8248
rect 419534 8236 419540 8248
rect 419592 8236 419598 8288
rect 74994 8168 75000 8220
rect 75052 8208 75058 8220
rect 423674 8208 423680 8220
rect 75052 8180 423680 8208
rect 75052 8168 75058 8180
rect 423674 8168 423680 8180
rect 423732 8168 423738 8220
rect 85666 8100 85672 8152
rect 85724 8140 85730 8152
rect 434714 8140 434720 8152
rect 85724 8112 434720 8140
rect 85724 8100 85730 8112
rect 434714 8100 434720 8112
rect 434772 8100 434778 8152
rect 82078 8032 82084 8084
rect 82136 8072 82142 8084
rect 430574 8072 430580 8084
rect 82136 8044 430580 8072
rect 82136 8032 82142 8044
rect 430574 8032 430580 8044
rect 430632 8032 430638 8084
rect 78582 7964 78588 8016
rect 78640 8004 78646 8016
rect 427814 8004 427820 8016
rect 78640 7976 427820 8004
rect 78640 7964 78646 7976
rect 427814 7964 427820 7976
rect 427872 7964 427878 8016
rect 92750 7896 92756 7948
rect 92808 7936 92814 7948
rect 442994 7936 443000 7948
rect 92808 7908 443000 7936
rect 92808 7896 92814 7908
rect 442994 7896 443000 7908
rect 443052 7896 443058 7948
rect 99834 7828 99840 7880
rect 99892 7868 99898 7880
rect 451274 7868 451280 7880
rect 99892 7840 451280 7868
rect 99892 7828 99898 7840
rect 451274 7828 451280 7840
rect 451332 7828 451338 7880
rect 114002 7760 114008 7812
rect 114060 7800 114066 7812
rect 466454 7800 466460 7812
rect 114060 7772 466460 7800
rect 114060 7760 114066 7772
rect 466454 7760 466460 7772
rect 466512 7760 466518 7812
rect 117590 7692 117596 7744
rect 117648 7732 117654 7744
rect 470594 7732 470600 7744
rect 117648 7704 470600 7732
rect 117648 7692 117654 7704
rect 470594 7692 470600 7704
rect 470652 7692 470658 7744
rect 106918 7624 106924 7676
rect 106976 7664 106982 7676
rect 459646 7664 459652 7676
rect 106976 7636 459652 7664
rect 106976 7624 106982 7636
rect 459646 7624 459652 7636
rect 459704 7624 459710 7676
rect 124674 7556 124680 7608
rect 124732 7596 124738 7608
rect 478874 7596 478880 7608
rect 124732 7568 478880 7596
rect 124732 7556 124738 7568
rect 478874 7556 478880 7568
rect 478932 7556 478938 7608
rect 64322 7488 64328 7540
rect 64380 7528 64386 7540
rect 411254 7528 411260 7540
rect 64380 7500 411260 7528
rect 64380 7488 64386 7500
rect 411254 7488 411260 7500
rect 411312 7488 411318 7540
rect 60826 7420 60832 7472
rect 60884 7460 60890 7472
rect 407114 7460 407120 7472
rect 60884 7432 407120 7460
rect 60884 7420 60890 7432
rect 407114 7420 407120 7432
rect 407172 7420 407178 7472
rect 50154 7352 50160 7404
rect 50212 7392 50218 7404
rect 396074 7392 396080 7404
rect 50212 7364 396080 7392
rect 50212 7352 50218 7364
rect 396074 7352 396080 7364
rect 396132 7352 396138 7404
rect 57238 7284 57244 7336
rect 57296 7324 57302 7336
rect 402974 7324 402980 7336
rect 57296 7296 402980 7324
rect 57296 7284 57302 7296
rect 402974 7284 402980 7296
rect 403032 7284 403038 7336
rect 43070 7216 43076 7268
rect 43128 7256 43134 7268
rect 387794 7256 387800 7268
rect 43128 7228 387800 7256
rect 43128 7216 43134 7228
rect 387794 7216 387800 7228
rect 387852 7216 387858 7268
rect 39574 7148 39580 7200
rect 39632 7188 39638 7200
rect 383654 7188 383660 7200
rect 39632 7160 383660 7188
rect 39632 7148 39638 7160
rect 383654 7148 383660 7160
rect 383712 7148 383718 7200
rect 41874 7080 41880 7132
rect 41932 7120 41938 7132
rect 386414 7120 386420 7132
rect 41932 7092 386420 7120
rect 41932 7080 41938 7092
rect 386414 7080 386420 7092
rect 386472 7080 386478 7132
rect 20622 7012 20628 7064
rect 20680 7052 20686 7064
rect 362954 7052 362960 7064
rect 20680 7024 362960 7052
rect 20680 7012 20686 7024
rect 362954 7012 362960 7024
rect 363012 7012 363018 7064
rect 73798 6808 73804 6860
rect 73856 6848 73862 6860
rect 422294 6848 422300 6860
rect 73856 6820 422300 6848
rect 73856 6808 73862 6820
rect 422294 6808 422300 6820
rect 422352 6808 422358 6860
rect 84470 6740 84476 6792
rect 84528 6780 84534 6792
rect 433334 6780 433340 6792
rect 84528 6752 433340 6780
rect 84528 6740 84534 6752
rect 433334 6740 433340 6752
rect 433392 6740 433398 6792
rect 77386 6672 77392 6724
rect 77444 6712 77450 6724
rect 426434 6712 426440 6724
rect 77444 6684 426440 6712
rect 77444 6672 77450 6684
rect 426434 6672 426440 6684
rect 426492 6672 426498 6724
rect 80882 6604 80888 6656
rect 80940 6644 80946 6656
rect 429286 6644 429292 6656
rect 80940 6616 429292 6644
rect 80940 6604 80946 6616
rect 429286 6604 429292 6616
rect 429344 6604 429350 6656
rect 91554 6536 91560 6588
rect 91612 6576 91618 6588
rect 441614 6576 441620 6588
rect 91612 6548 441620 6576
rect 91612 6536 91618 6548
rect 441614 6536 441620 6548
rect 441672 6536 441678 6588
rect 87966 6468 87972 6520
rect 88024 6508 88030 6520
rect 437474 6508 437480 6520
rect 88024 6480 437480 6508
rect 88024 6468 88030 6480
rect 437474 6468 437480 6480
rect 437532 6468 437538 6520
rect 98638 6400 98644 6452
rect 98696 6440 98702 6452
rect 449894 6440 449900 6452
rect 98696 6412 449900 6440
rect 98696 6400 98702 6412
rect 449894 6400 449900 6412
rect 449952 6400 449958 6452
rect 109310 6332 109316 6384
rect 109368 6372 109374 6384
rect 460934 6372 460940 6384
rect 109368 6344 460940 6372
rect 109368 6332 109374 6344
rect 460934 6332 460940 6344
rect 460992 6332 460998 6384
rect 95142 6264 95148 6316
rect 95200 6304 95206 6316
rect 445754 6304 445760 6316
rect 95200 6276 445760 6304
rect 95200 6264 95206 6276
rect 445754 6264 445760 6276
rect 445812 6264 445818 6316
rect 102226 6196 102232 6248
rect 102284 6236 102290 6248
rect 454034 6236 454040 6248
rect 102284 6208 454040 6236
rect 102284 6196 102290 6208
rect 454034 6196 454040 6208
rect 454092 6196 454098 6248
rect 116394 6128 116400 6180
rect 116452 6168 116458 6180
rect 469214 6168 469220 6180
rect 116452 6140 469220 6168
rect 116452 6128 116458 6140
rect 469214 6128 469220 6140
rect 469272 6128 469278 6180
rect 70302 6060 70308 6112
rect 70360 6100 70366 6112
rect 418154 6100 418160 6112
rect 70360 6072 418160 6100
rect 70360 6060 70366 6072
rect 418154 6060 418160 6072
rect 418212 6060 418218 6112
rect 63218 5992 63224 6044
rect 63276 6032 63282 6044
rect 409874 6032 409880 6044
rect 63276 6004 409880 6032
rect 63276 5992 63282 6004
rect 409874 5992 409880 6004
rect 409932 5992 409938 6044
rect 66714 5924 66720 5976
rect 66772 5964 66778 5976
rect 414014 5964 414020 5976
rect 66772 5936 414020 5964
rect 66772 5924 66778 5936
rect 414014 5924 414020 5936
rect 414072 5924 414078 5976
rect 48958 5856 48964 5908
rect 49016 5896 49022 5908
rect 394694 5896 394700 5908
rect 49016 5868 394700 5896
rect 49016 5856 49022 5868
rect 394694 5856 394700 5868
rect 394752 5856 394758 5908
rect 59630 5788 59636 5840
rect 59688 5828 59694 5840
rect 405734 5828 405740 5840
rect 59688 5800 405740 5828
rect 59688 5788 59694 5800
rect 405734 5788 405740 5800
rect 405792 5788 405798 5840
rect 56042 5720 56048 5772
rect 56100 5760 56106 5772
rect 401594 5760 401600 5772
rect 56100 5732 401600 5760
rect 56100 5720 56106 5732
rect 401594 5720 401600 5732
rect 401652 5720 401658 5772
rect 52546 5652 52552 5704
rect 52604 5692 52610 5704
rect 397546 5692 397552 5704
rect 52604 5664 397552 5692
rect 52604 5652 52610 5664
rect 397546 5652 397552 5664
rect 397604 5652 397610 5704
rect 13538 5584 13544 5636
rect 13596 5624 13602 5636
rect 354674 5624 354680 5636
rect 13596 5596 354680 5624
rect 13596 5584 13602 5596
rect 354674 5584 354680 5596
rect 354732 5584 354738 5636
rect 90358 5448 90364 5500
rect 90416 5488 90422 5500
rect 440234 5488 440240 5500
rect 90416 5460 440240 5488
rect 90416 5448 90422 5460
rect 440234 5448 440240 5460
rect 440292 5448 440298 5500
rect 86862 5380 86868 5432
rect 86920 5420 86926 5432
rect 436094 5420 436100 5432
rect 86920 5392 436100 5420
rect 86920 5380 86926 5392
rect 436094 5380 436100 5392
rect 436152 5380 436158 5432
rect 79686 5312 79692 5364
rect 79744 5352 79750 5364
rect 429194 5352 429200 5364
rect 79744 5324 429200 5352
rect 79744 5312 79750 5324
rect 429194 5312 429200 5324
rect 429252 5312 429258 5364
rect 101030 5244 101036 5296
rect 101088 5284 101094 5296
rect 452654 5284 452660 5296
rect 101088 5256 452660 5284
rect 101088 5244 101094 5256
rect 452654 5244 452660 5256
rect 452712 5244 452718 5296
rect 108114 5176 108120 5228
rect 108172 5216 108178 5228
rect 459554 5216 459560 5228
rect 108172 5188 459560 5216
rect 108172 5176 108178 5188
rect 459554 5176 459560 5188
rect 459612 5176 459618 5228
rect 97442 5108 97448 5160
rect 97500 5148 97506 5160
rect 448514 5148 448520 5160
rect 97500 5120 448520 5148
rect 97500 5108 97506 5120
rect 448514 5108 448520 5120
rect 448572 5108 448578 5160
rect 118786 5040 118792 5092
rect 118844 5080 118850 5092
rect 471974 5080 471980 5092
rect 118844 5052 471980 5080
rect 118844 5040 118850 5052
rect 471974 5040 471980 5052
rect 472032 5040 472038 5092
rect 115198 4972 115204 5024
rect 115256 5012 115262 5024
rect 467834 5012 467840 5024
rect 115256 4984 467840 5012
rect 115256 4972 115262 4984
rect 467834 4972 467840 4984
rect 467892 4972 467898 5024
rect 111610 4904 111616 4956
rect 111668 4944 111674 4956
rect 463694 4944 463700 4956
rect 111668 4916 463700 4944
rect 111668 4904 111674 4916
rect 463694 4904 463700 4916
rect 463752 4904 463758 4956
rect 104526 4836 104532 4888
rect 104584 4876 104590 4888
rect 456794 4876 456800 4888
rect 104584 4848 456800 4876
rect 104584 4836 104590 4848
rect 456794 4836 456800 4848
rect 456852 4836 456858 4888
rect 122282 4768 122288 4820
rect 122340 4808 122346 4820
rect 476114 4808 476120 4820
rect 122340 4780 476120 4808
rect 122340 4768 122346 4780
rect 476114 4768 476120 4780
rect 476172 4768 476178 4820
rect 93946 4700 93952 4752
rect 94004 4740 94010 4752
rect 444374 4740 444380 4752
rect 94004 4712 444380 4740
rect 94004 4700 94010 4712
rect 444374 4700 444380 4712
rect 444432 4700 444438 4752
rect 83274 4632 83280 4684
rect 83332 4672 83338 4684
rect 431954 4672 431960 4684
rect 83332 4644 431960 4672
rect 83332 4632 83338 4644
rect 431954 4632 431960 4644
rect 432012 4632 432018 4684
rect 76190 4564 76196 4616
rect 76248 4604 76254 4616
rect 425054 4604 425060 4616
rect 76248 4576 425060 4604
rect 76248 4564 76254 4576
rect 425054 4564 425060 4576
rect 425112 4564 425118 4616
rect 72602 4496 72608 4548
rect 72660 4536 72666 4548
rect 420914 4536 420920 4548
rect 72660 4508 420920 4536
rect 72660 4496 72666 4508
rect 420914 4496 420920 4508
rect 420972 4496 420978 4548
rect 69106 4428 69112 4480
rect 69164 4468 69170 4480
rect 416774 4468 416780 4480
rect 69164 4440 416780 4468
rect 69164 4428 69170 4440
rect 416774 4428 416780 4440
rect 416832 4428 416838 4480
rect 21818 4360 21824 4412
rect 21876 4400 21882 4412
rect 364334 4400 364340 4412
rect 21876 4372 364340 4400
rect 21876 4360 21882 4372
rect 364334 4360 364340 4372
rect 364392 4360 364398 4412
rect 12342 4292 12348 4344
rect 12400 4332 12406 4344
rect 353294 4332 353300 4344
rect 12400 4304 353300 4332
rect 12400 4292 12406 4304
rect 353294 4292 353300 4304
rect 353352 4292 353358 4344
rect 17034 4224 17040 4276
rect 17092 4264 17098 4276
rect 358814 4264 358820 4276
rect 17092 4236 358820 4264
rect 17092 4224 17098 4236
rect 358814 4224 358820 4236
rect 358872 4224 358878 4276
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 7558 4128 7564 4140
rect 1728 4100 7564 4128
rect 1728 4088 1734 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 351914 4128 351920 4140
rect 11204 4100 351920 4128
rect 11204 4088 11210 4100
rect 351914 4088 351920 4100
rect 351972 4088 351978 4140
rect 26510 4020 26516 4072
rect 26568 4060 26574 4072
rect 27522 4060 27528 4072
rect 26568 4032 27528 4060
rect 26568 4020 26574 4032
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 27617 4063 27675 4069
rect 27617 4029 27629 4063
rect 27663 4060 27675 4063
rect 367186 4060 367192 4072
rect 27663 4032 367192 4060
rect 27663 4029 27675 4032
rect 27617 4023 27675 4029
rect 367186 4020 367192 4032
rect 367244 4020 367250 4072
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 357434 3992 357440 4004
rect 15988 3964 357440 3992
rect 15988 3952 15994 3964
rect 357434 3952 357440 3964
rect 357492 3952 357498 4004
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 356054 3924 356060 3936
rect 14792 3896 356060 3924
rect 14792 3884 14798 3896
rect 356054 3884 356060 3896
rect 356112 3884 356118 3936
rect 25314 3816 25320 3868
rect 25372 3856 25378 3868
rect 27617 3859 27675 3865
rect 27617 3856 27629 3859
rect 25372 3828 27629 3856
rect 25372 3816 25378 3828
rect 27617 3825 27629 3828
rect 27663 3825 27675 3859
rect 27617 3819 27675 3825
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 371234 3856 371240 3868
rect 28960 3828 371240 3856
rect 28960 3816 28966 3828
rect 371234 3816 371240 3828
rect 371292 3816 371298 3868
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 375374 3788 375380 3800
rect 32456 3760 375380 3788
rect 32456 3748 32462 3760
rect 375374 3748 375380 3760
rect 375432 3748 375438 3800
rect 105722 3680 105728 3732
rect 105780 3720 105786 3732
rect 106182 3720 106188 3732
rect 105780 3692 106188 3720
rect 105780 3680 105786 3692
rect 106182 3680 106188 3692
rect 106240 3680 106246 3732
rect 123478 3680 123484 3732
rect 123536 3720 123542 3732
rect 124122 3720 124128 3732
rect 123536 3692 124128 3720
rect 123536 3680 123542 3692
rect 124122 3680 124128 3692
rect 124180 3680 124186 3732
rect 125137 3723 125195 3729
rect 125137 3689 125149 3723
rect 125183 3720 125195 3723
rect 465718 3720 465724 3732
rect 125183 3692 465724 3720
rect 125183 3689 125195 3692
rect 125137 3683 125195 3689
rect 465718 3680 465724 3692
rect 465776 3680 465782 3732
rect 53742 3612 53748 3664
rect 53800 3652 53806 3664
rect 398834 3652 398840 3664
rect 53800 3624 398840 3652
rect 53800 3612 53806 3624
rect 398834 3612 398840 3624
rect 398892 3612 398898 3664
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 18598 3584 18604 3596
rect 8812 3556 18604 3584
rect 8812 3544 8818 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 39298 3584 39304 3596
rect 34848 3556 39304 3584
rect 34848 3544 34854 3556
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 46658 3544 46664 3596
rect 46716 3584 46722 3596
rect 391934 3584 391940 3596
rect 46716 3556 391940 3584
rect 46716 3544 46722 3556
rect 391934 3544 391940 3556
rect 391992 3544 391998 3596
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 14458 3516 14464 3528
rect 2924 3488 14464 3516
rect 2924 3476 2930 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 22738 3516 22744 3528
rect 18288 3488 22744 3516
rect 18288 3476 18294 3488
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 32306 3516 32312 3528
rect 27764 3488 32312 3516
rect 27764 3476 27770 3488
rect 32306 3476 32312 3488
rect 32364 3476 32370 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 438854 3516 438860 3528
rect 89220 3488 438860 3516
rect 89220 3476 89226 3488
rect 438854 3476 438860 3488
rect 438912 3476 438918 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 17218 3448 17224 3460
rect 624 3420 17224 3448
rect 624 3408 630 3420
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 35158 3448 35164 3460
rect 31352 3420 35164 3448
rect 31352 3408 31358 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 43438 3448 43444 3460
rect 38436 3420 43444 3448
rect 38436 3408 38442 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 96246 3408 96252 3460
rect 96304 3448 96310 3460
rect 447134 3448 447140 3460
rect 96304 3420 447140 3448
rect 96304 3408 96310 3420
rect 447134 3408 447140 3420
rect 447192 3408 447198 3460
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 338850 3380 338856 3392
rect 6512 3352 338856 3380
rect 6512 3340 6518 3352
rect 338850 3340 338856 3352
rect 338908 3340 338914 3392
rect 5258 3272 5264 3324
rect 5316 3312 5322 3324
rect 336090 3312 336096 3324
rect 5316 3284 336096 3312
rect 5316 3272 5322 3284
rect 336090 3272 336096 3284
rect 336148 3272 336154 3324
rect 327718 3244 327724 3256
rect 22066 3216 327724 3244
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 22066 3108 22094 3216
rect 327718 3204 327724 3216
rect 327776 3204 327782 3256
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 331858 3176 331864 3188
rect 24268 3148 331864 3176
rect 24268 3136 24274 3148
rect 331858 3136 331864 3148
rect 331916 3136 331922 3188
rect 19484 3080 22094 3108
rect 19484 3068 19490 3080
rect 35986 3068 35992 3120
rect 36044 3108 36050 3120
rect 334618 3108 334624 3120
rect 36044 3080 334624 3108
rect 36044 3068 36050 3080
rect 334618 3068 334624 3080
rect 334676 3068 334682 3120
rect 67910 3000 67916 3052
rect 67968 3040 67974 3052
rect 322290 3040 322296 3052
rect 67968 3012 322296 3040
rect 67968 3000 67974 3012
rect 322290 3000 322296 3012
rect 322348 3000 322354 3052
rect 103330 2932 103336 2984
rect 103388 2972 103394 2984
rect 323670 2972 323676 2984
rect 103388 2944 323676 2972
rect 103388 2932 103394 2944
rect 323670 2932 323676 2944
rect 323728 2932 323734 2984
rect 110506 2864 110512 2916
rect 110564 2904 110570 2916
rect 324958 2904 324964 2916
rect 110564 2876 324964 2904
rect 110564 2864 110570 2876
rect 324958 2864 324964 2876
rect 325016 2864 325022 2916
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 125137 2839 125195 2845
rect 125137 2836 125149 2839
rect 121144 2808 125149 2836
rect 121144 2796 121150 2808
rect 125137 2805 125149 2808
rect 125183 2805 125195 2839
rect 125137 2799 125195 2805
<< via1 >>
rect 332508 700952 332560 701004
rect 472072 700952 472124 701004
rect 283840 700884 283892 700936
rect 469220 700884 469272 700936
rect 267648 700816 267700 700868
rect 470600 700816 470652 700868
rect 218980 700748 219032 700800
rect 467932 700748 467984 700800
rect 202788 700680 202840 700732
rect 467840 700680 467892 700732
rect 154120 700612 154172 700664
rect 465080 700612 465132 700664
rect 56784 700544 56836 700596
rect 105544 700544 105596 700596
rect 137836 700544 137888 700596
rect 466460 700544 466512 700596
rect 89168 700476 89220 700528
rect 462228 700476 462280 700528
rect 72976 700408 73028 700460
rect 463700 700408 463752 700460
rect 24308 700340 24360 700392
rect 460940 700340 460992 700392
rect 8116 700272 8168 700324
rect 462412 700340 462464 700392
rect 462320 700272 462372 700324
rect 472808 700272 472860 700324
rect 530584 700272 530636 700324
rect 543464 700272 543516 700324
rect 348792 700204 348844 700256
rect 471980 700204 472032 700256
rect 397460 700136 397512 700188
rect 472716 700136 472768 700188
rect 413652 700068 413704 700120
rect 472900 700068 472952 700120
rect 446128 700000 446180 700052
rect 491300 700000 491352 700052
rect 250444 699660 250496 699712
rect 251456 699660 251508 699712
rect 475384 699660 475436 699712
rect 478512 699660 478564 699712
rect 527180 699660 527232 699712
rect 528560 699660 528612 699712
rect 536104 696940 536156 696992
rect 580172 696940 580224 696992
rect 529204 683136 529256 683188
rect 580172 683136 580224 683188
rect 276296 682388 276348 682440
rect 316040 682388 316092 682440
rect 267188 681708 267240 681760
rect 276296 681708 276348 681760
rect 276756 681708 276808 681760
rect 455328 680348 455380 680400
rect 483480 680348 483532 680400
rect 97908 679260 97960 679312
rect 99656 679260 99708 679312
rect 241428 679260 241480 679312
rect 316684 679260 316736 679312
rect 85488 678988 85540 679040
rect 316776 678988 316828 679040
rect 88064 677288 88116 677340
rect 93860 677288 93912 677340
rect 271880 676268 271932 676320
rect 272892 676268 272944 676320
rect 78588 675452 78640 675504
rect 86132 675452 86184 675504
rect 238668 675452 238720 675504
rect 241520 675452 241572 675504
rect 505560 674296 505612 674348
rect 506388 674296 506440 674348
rect 482928 674160 482980 674212
rect 490656 674160 490708 674212
rect 477408 674092 477460 674144
rect 487252 674092 487304 674144
rect 493324 673888 493376 673940
rect 494428 673888 494480 673940
rect 499488 673480 499540 673532
rect 500224 673480 500276 673532
rect 82728 672732 82780 672784
rect 90640 672732 90692 672784
rect 92388 672732 92440 672784
rect 96712 672732 96764 672784
rect 114744 672528 114796 672580
rect 115848 672528 115900 672580
rect 242808 672052 242860 672104
rect 246304 672052 246356 672104
rect 251180 672052 251232 672104
rect 252192 672052 252244 672104
rect 258540 672052 258592 672104
rect 259368 672052 259420 672104
rect 3516 670692 3568 670744
rect 323676 670692 323728 670744
rect 3424 656888 3476 656940
rect 336096 656888 336148 656940
rect 533344 643084 533396 643136
rect 580172 643084 580224 643136
rect 502248 632884 502300 632936
rect 511448 632884 511500 632936
rect 264888 632816 264940 632868
rect 272064 632816 272116 632868
rect 502432 632816 502484 632868
rect 516324 632816 516376 632868
rect 270408 632748 270460 632800
rect 281540 632748 281592 632800
rect 506388 632748 506440 632800
rect 521292 632748 521344 632800
rect 111892 632680 111944 632732
rect 116584 632680 116636 632732
rect 117688 632680 117740 632732
rect 126428 632680 126480 632732
rect 271972 632680 272024 632732
rect 286324 632680 286376 632732
rect 506480 632680 506532 632732
rect 526168 632680 526220 632732
rect 486884 632340 486936 632392
rect 491576 632340 491628 632392
rect 247684 632272 247736 632324
rect 248420 632272 248472 632324
rect 260840 632136 260892 632188
rect 266728 632136 266780 632188
rect 499580 632136 499632 632188
rect 506572 632136 506624 632188
rect 78036 632068 78088 632120
rect 78588 632068 78640 632120
rect 108948 632068 109000 632120
rect 111800 632068 111852 632120
rect 115848 632068 115900 632120
rect 121552 632068 121604 632120
rect 237932 632068 237984 632120
rect 238668 632068 238720 632120
rect 255320 632068 255372 632120
rect 256884 632068 256936 632120
rect 259368 632068 259420 632120
rect 261760 632068 261812 632120
rect 482008 632068 482060 632120
rect 482928 632068 482980 632120
rect 491852 632068 491904 632120
rect 493324 632068 493376 632120
rect 500224 632068 500276 632120
rect 501604 632068 501656 632120
rect 538864 630640 538916 630692
rect 580172 630640 580224 630692
rect 72792 628260 72844 628312
rect 232872 628260 232924 628312
rect 72700 628192 72752 628244
rect 130384 628192 130436 628244
rect 232688 628192 232740 628244
rect 289268 628192 289320 628244
rect 73068 628124 73120 628176
rect 130568 628124 130620 628176
rect 233148 628124 233200 628176
rect 290372 628124 290424 628176
rect 72608 628056 72660 628108
rect 133144 628056 133196 628108
rect 235264 628056 235316 628108
rect 290464 628056 290516 628108
rect 74448 627988 74500 628040
rect 232872 627988 232924 628040
rect 313924 627988 313976 628040
rect 232780 627920 232832 627972
rect 320824 627920 320876 627972
rect 233148 627852 233200 627904
rect 72976 627648 73028 627700
rect 129004 627648 129056 627700
rect 233056 627648 233108 627700
rect 289084 627648 289136 627700
rect 72884 627580 72936 627632
rect 130476 627580 130528 627632
rect 232964 627580 233016 627632
rect 289176 627580 289228 627632
rect 290464 627172 290516 627224
rect 454040 627172 454092 627224
rect 454040 626560 454092 626612
rect 472624 626560 472676 626612
rect 133144 623704 133196 623756
rect 232780 623704 232832 623756
rect 320824 623024 320876 623076
rect 472164 623024 472216 623076
rect 472532 623024 472584 623076
rect 130568 619556 130620 619608
rect 232320 619556 232372 619608
rect 289268 618876 289320 618928
rect 451280 618876 451332 618928
rect 452200 618876 452252 618928
rect 452200 618264 452252 618316
rect 472624 618264 472676 618316
rect 313924 614728 313976 614780
rect 472256 614728 472308 614780
rect 472532 614728 472584 614780
rect 130476 611260 130528 611312
rect 232964 611260 233016 611312
rect 289176 610580 289228 610632
rect 449900 610580 449952 610632
rect 449900 609968 449952 610020
rect 472624 609968 472676 610020
rect 129004 607112 129056 607164
rect 232412 607112 232464 607164
rect 289084 606432 289136 606484
rect 472440 606432 472492 606484
rect 130384 603032 130436 603084
rect 233148 603032 233200 603084
rect 290464 602352 290516 602404
rect 447140 602352 447192 602404
rect 447140 601672 447192 601724
rect 472624 601672 472676 601724
rect 445024 589296 445076 589348
rect 472624 589296 472676 589348
rect 459468 585148 459520 585200
rect 472624 585148 472676 585200
rect 72792 582224 72844 582276
rect 72976 582224 73028 582276
rect 444380 578144 444432 578196
rect 445024 578144 445076 578196
rect 472532 578144 472584 578196
rect 472992 578144 473044 578196
rect 472440 578076 472492 578128
rect 473084 578076 473136 578128
rect 231768 577736 231820 577788
rect 472532 577804 472584 577856
rect 72884 577668 72936 577720
rect 232964 577668 233016 577720
rect 72976 577600 73028 577652
rect 232780 577600 232832 577652
rect 444380 577600 444432 577652
rect 72792 577532 72844 577584
rect 231768 577532 231820 577584
rect 472440 577532 472492 577584
rect 75828 577464 75880 577516
rect 233148 577464 233200 577516
rect 235264 577464 235316 577516
rect 472624 577464 472676 577516
rect 73068 577396 73120 577448
rect 233056 577396 233108 577448
rect 17868 576852 17920 576904
rect 71780 576852 71832 576904
rect 537484 576852 537536 576904
rect 580172 576852 580224 576904
rect 233056 576172 233108 576224
rect 339408 576172 339460 576224
rect 3516 576104 3568 576156
rect 331864 576104 331916 576156
rect 475384 576104 475436 576156
rect 480168 576104 480220 576156
rect 528560 576104 528612 576156
rect 475384 575832 475436 575884
rect 339408 575424 339460 575476
rect 473176 575424 473228 575476
rect 86132 573996 86184 574048
rect 360292 573996 360344 574048
rect 426348 573996 426400 574048
rect 519636 573996 519688 574048
rect 76380 573928 76432 573980
rect 351920 573928 351972 573980
rect 367008 573928 367060 573980
rect 488540 573928 488592 573980
rect 89444 573860 89496 573912
rect 367100 573860 367152 573912
rect 369768 573860 369820 573912
rect 490196 573860 490248 573912
rect 114008 573792 114060 573844
rect 395344 573792 395396 573844
rect 407028 573792 407080 573844
rect 509792 573792 509844 573844
rect 112352 573724 112404 573776
rect 399484 573724 399536 573776
rect 404268 573724 404320 573776
rect 508136 573724 508188 573776
rect 120540 573656 120592 573708
rect 410524 573656 410576 573708
rect 416688 573656 416740 573708
rect 514668 573656 514720 573708
rect 117228 573588 117280 573640
rect 407764 573588 407816 573640
rect 411904 573588 411956 573640
rect 511448 573588 511500 573640
rect 122196 573520 122248 573572
rect 417424 573520 417476 573572
rect 419448 573520 419500 573572
rect 516324 573520 516376 573572
rect 118516 573452 118568 573504
rect 413284 573452 413336 573504
rect 414664 573452 414716 573504
rect 513104 573452 513156 573504
rect 123760 573384 123812 573436
rect 421564 573384 421616 573436
rect 423588 573384 423640 573436
rect 517980 573384 518032 573436
rect 125416 573316 125468 573368
rect 431224 573316 431276 573368
rect 433248 573316 433300 573368
rect 522856 573316 522908 573368
rect 84108 573248 84160 573300
rect 357440 573248 357492 573300
rect 429108 573248 429160 573300
rect 521292 573248 521344 573300
rect 87788 573180 87840 573232
rect 104164 573180 104216 573232
rect 106924 573180 106976 573232
rect 115572 573180 115624 573232
rect 363604 573180 363656 573232
rect 436008 573180 436060 573232
rect 524512 573180 524564 573232
rect 82728 573112 82780 573164
rect 327724 573112 327776 573164
rect 438768 573112 438820 573164
rect 526168 573112 526220 573164
rect 331956 573044 332008 573096
rect 441528 573044 441580 573096
rect 527824 573044 527876 573096
rect 91008 572976 91060 573028
rect 334716 572976 334768 573028
rect 409144 572976 409196 573028
rect 478696 572976 478748 573028
rect 482284 572976 482336 573028
rect 491760 572976 491812 573028
rect 81256 572908 81308 572960
rect 322204 572908 322256 572960
rect 420184 572908 420236 572960
rect 480352 572908 480404 572960
rect 485228 572908 485280 572960
rect 102508 572840 102560 572892
rect 105544 572840 105596 572892
rect 126888 572840 126940 572892
rect 323584 572840 323636 572892
rect 443644 572840 443696 572892
rect 482008 572840 482060 572892
rect 100668 572772 100720 572824
rect 104164 572772 104216 572824
rect 128728 572772 128780 572824
rect 324964 572772 325016 572824
rect 476764 572772 476816 572824
rect 483572 572772 483624 572824
rect 77944 572704 77996 572756
rect 78588 572704 78640 572756
rect 94320 572704 94372 572756
rect 95148 572704 95200 572756
rect 95976 572704 96028 572756
rect 97264 572704 97316 572756
rect 97632 572704 97684 572756
rect 98644 572704 98696 572756
rect 99288 572704 99340 572756
rect 101404 572704 101456 572756
rect 105820 572704 105872 572756
rect 108304 572704 108356 572756
rect 108948 572704 109000 572756
rect 111064 572704 111116 572756
rect 237840 572704 237892 572756
rect 238668 572704 238720 572756
rect 246028 572704 246080 572756
rect 246948 572704 247000 572756
rect 255872 572704 255924 572756
rect 256608 572704 256660 572756
rect 264060 572704 264112 572756
rect 264888 572704 264940 572756
rect 272248 572704 272300 572756
rect 273168 572704 273220 572756
rect 273904 572704 273956 572756
rect 274548 572704 274600 572756
rect 275468 572704 275520 572756
rect 275928 572704 275980 572756
rect 280436 572704 280488 572756
rect 281448 572704 281500 572756
rect 282092 572704 282144 572756
rect 282828 572704 282880 572756
rect 283656 572704 283708 572756
rect 284208 572704 284260 572756
rect 478144 572704 478196 572756
rect 480904 572704 480956 572756
rect 486884 572704 486936 572756
rect 497464 572704 497516 572756
rect 498384 572704 498436 572756
rect 247684 572636 247736 572688
rect 349804 572636 349856 572688
rect 236276 572568 236328 572620
rect 341524 572568 341576 572620
rect 239496 572500 239548 572552
rect 345020 572500 345072 572552
rect 244188 572432 244240 572484
rect 356060 572432 356112 572484
rect 257528 572364 257580 572416
rect 370504 572364 370556 572416
rect 382188 572364 382240 572416
rect 496728 572364 496780 572416
rect 254216 572296 254268 572348
rect 374644 572296 374696 572348
rect 379428 572296 379480 572348
rect 495072 572296 495124 572348
rect 262128 572228 262180 572280
rect 388444 572228 388496 572280
rect 265716 572160 265768 572212
rect 396724 572160 396776 572212
rect 340788 572092 340840 572144
rect 477040 572092 477092 572144
rect 110328 572024 110380 572076
rect 382924 572024 382976 572076
rect 107384 571956 107436 572008
rect 393964 571956 394016 572008
rect 3240 565836 3292 565888
rect 334624 565836 334676 565888
rect 3332 553392 3384 553444
rect 322296 553392 322348 553444
rect 482376 536800 482428 536852
rect 579896 536800 579948 536852
rect 482468 524424 482520 524476
rect 580172 524424 580224 524476
rect 3516 500964 3568 501016
rect 320916 500964 320968 501016
rect 482560 484372 482612 484424
rect 580172 484372 580224 484424
rect 482652 470568 482704 470620
rect 580172 470568 580224 470620
rect 3516 462340 3568 462392
rect 330576 462340 330628 462392
rect 246948 456152 247000 456204
rect 353944 456152 353996 456204
rect 260748 456084 260800 456136
rect 387800 456084 387852 456136
rect 267648 456016 267700 456068
rect 400220 456016 400272 456068
rect 238668 453364 238720 453416
rect 340880 453364 340932 453416
rect 79968 453296 80020 453348
rect 342904 453296 342956 453348
rect 3516 448536 3568 448588
rect 325332 448536 325384 448588
rect 482744 430584 482796 430636
rect 579896 430584 579948 430636
rect 482836 418140 482888 418192
rect 580172 418140 580224 418192
rect 104164 412156 104216 412208
rect 389456 412156 389508 412208
rect 105544 412088 105596 412140
rect 392676 412088 392728 412140
rect 106924 412020 106976 412072
rect 396080 412020 396132 412072
rect 108304 411952 108356 412004
rect 398932 411952 398984 412004
rect 111064 411884 111116 411936
rect 405740 411884 405792 411936
rect 251088 411204 251140 411256
rect 369952 411204 370004 411256
rect 252468 411136 252520 411188
rect 371884 411136 371936 411188
rect 256608 411068 256660 411120
rect 378968 411068 379020 411120
rect 259368 411000 259420 411052
rect 385316 411000 385368 411052
rect 264888 410932 264940 410984
rect 394792 410932 394844 410984
rect 269028 410864 269080 410916
rect 403624 410864 403676 410916
rect 273168 410796 273220 410848
rect 410432 410796 410484 410848
rect 270408 410728 270460 410780
rect 407396 410728 407448 410780
rect 274548 410660 274600 410712
rect 414112 410660 414164 410712
rect 98644 410592 98696 410644
rect 383660 410592 383712 410644
rect 101404 410524 101456 410576
rect 386420 410524 386472 410576
rect 249708 410456 249760 410508
rect 364984 410456 365036 410508
rect 228824 410184 228876 410236
rect 327908 410184 327960 410236
rect 226248 410116 226300 410168
rect 326344 410116 326396 410168
rect 222108 410048 222160 410100
rect 325148 410048 325200 410100
rect 223488 409980 223540 410032
rect 329196 409980 329248 410032
rect 218980 409912 219032 409964
rect 332048 409912 332100 409964
rect 3148 409844 3200 409896
rect 329564 409844 329616 409896
rect 211068 409776 211120 409828
rect 333244 409776 333296 409828
rect 3700 409708 3752 409760
rect 328276 409708 328328 409760
rect 264888 409640 264940 409692
rect 319536 409640 319588 409692
rect 278688 409572 278740 409624
rect 337568 409572 337620 409624
rect 274548 409504 274600 409556
rect 336556 409504 336608 409556
rect 271788 409436 271840 409488
rect 335268 409436 335320 409488
rect 232872 409368 232924 409420
rect 459008 409368 459060 409420
rect 78588 409300 78640 409352
rect 342260 409300 342312 409352
rect 95148 409232 95200 409284
rect 376852 409232 376904 409284
rect 92388 409164 92440 409216
rect 374000 409164 374052 409216
rect 97264 409096 97316 409148
rect 379980 409096 380032 409148
rect 259368 409028 259420 409080
rect 326528 409028 326580 409080
rect 256608 408960 256660 409012
rect 324044 408960 324096 409012
rect 266268 408892 266320 408944
rect 337476 408892 337528 408944
rect 253848 408824 253900 408876
rect 330760 408824 330812 408876
rect 251088 408756 251140 408808
rect 329288 408756 329340 408808
rect 213828 408688 213880 408740
rect 321008 408688 321060 408740
rect 216588 408620 216640 408672
rect 337384 408620 337436 408672
rect 286508 408552 286560 408604
rect 319444 408552 319496 408604
rect 276848 408484 276900 408536
rect 322572 408484 322624 408536
rect 114468 408416 114520 408468
rect 332416 408416 332468 408468
rect 124128 408348 124180 408400
rect 318248 408348 318300 408400
rect 284208 408280 284260 408332
rect 328000 408280 328052 408332
rect 269028 408212 269080 408264
rect 318432 408212 318484 408264
rect 262128 408144 262180 408196
rect 319628 408144 319680 408196
rect 249708 408076 249760 408128
rect 325424 408076 325476 408128
rect 246948 408008 247000 408060
rect 336280 408008 336332 408060
rect 140688 407940 140740 407992
rect 157524 407940 157576 407992
rect 234528 407940 234580 407992
rect 323860 407940 323912 407992
rect 139308 407872 139360 407924
rect 157432 407872 157484 407924
rect 241428 407872 241480 407924
rect 332232 407872 332284 407924
rect 71688 407804 71740 407856
rect 156788 407804 156840 407856
rect 237288 407804 237340 407856
rect 334900 407804 334952 407856
rect 66168 407736 66220 407788
rect 156696 407736 156748 407788
rect 231768 407736 231820 407788
rect 330852 407736 330904 407788
rect 64512 407668 64564 407720
rect 156604 407668 156656 407720
rect 209504 407668 209556 407720
rect 327816 407668 327868 407720
rect 121368 407600 121420 407652
rect 322664 407600 322716 407652
rect 117228 407532 117280 407584
rect 318524 407532 318576 407584
rect 126888 407464 126940 407516
rect 329472 407464 329524 407516
rect 118608 407396 118660 407448
rect 321376 407396 321428 407448
rect 111708 407328 111760 407380
rect 328184 407328 328236 407380
rect 108948 407260 109000 407312
rect 325516 407260 325568 407312
rect 300768 407192 300820 407244
rect 317604 407192 317656 407244
rect 151360 407124 151412 407176
rect 161480 407124 161532 407176
rect 299388 407124 299440 407176
rect 317512 407124 317564 407176
rect 52368 407056 52420 407108
rect 166264 407056 166316 407108
rect 282828 407056 282880 407108
rect 429476 407056 429528 407108
rect 56508 406988 56560 407040
rect 170404 406988 170456 407040
rect 284116 406988 284168 407040
rect 432696 406988 432748 407040
rect 59268 406920 59320 406972
rect 173164 406920 173216 406972
rect 285588 406920 285640 406972
rect 436192 406920 436244 406972
rect 53472 406852 53524 406904
rect 169024 406852 169076 406904
rect 286968 406852 287020 406904
rect 438952 406852 439004 406904
rect 61108 406784 61160 406836
rect 178408 406784 178460 406836
rect 288348 406784 288400 406836
rect 442172 406784 442224 406836
rect 99288 406716 99340 406768
rect 332324 406716 332376 406768
rect 95976 406648 96028 406700
rect 334992 406648 335044 406700
rect 86224 406580 86276 406632
rect 326436 406580 326488 406632
rect 83648 406512 83700 406564
rect 323952 406512 324004 406564
rect 88616 406444 88668 406496
rect 336188 406444 336240 406496
rect 81072 406376 81124 406428
rect 332140 406376 332192 406428
rect 48688 406308 48740 406360
rect 162124 406308 162176 406360
rect 281448 406308 281500 406360
rect 426440 406308 426492 406360
rect 278596 406240 278648 406292
rect 423772 406240 423824 406292
rect 277308 406172 277360 406224
rect 420000 406172 420052 406224
rect 275928 406104 275980 406156
rect 416872 406104 416924 406156
rect 242808 406036 242860 406088
rect 353668 406036 353720 406088
rect 241336 405968 241388 406020
rect 349436 405968 349488 406020
rect 238576 405900 238628 405952
rect 322388 405900 322440 405952
rect 243728 405832 243780 405884
rect 321284 405832 321336 405884
rect 281080 405764 281132 405816
rect 318340 405764 318392 405816
rect 397368 403656 397420 403708
rect 503720 403656 503772 403708
rect 394424 403588 394476 403640
rect 502340 403588 502392 403640
rect 400772 402500 400824 402552
rect 506480 402500 506532 402552
rect 391296 402432 391348 402484
rect 500960 402432 501012 402484
rect 388076 402364 388128 402416
rect 499580 402364 499632 402416
rect 384948 402296 385000 402348
rect 497464 402296 497516 402348
rect 375288 402228 375340 402280
rect 492680 402228 492732 402280
rect 320088 401616 320140 401668
rect 323768 401616 323820 401668
rect 349068 401548 349120 401600
rect 420184 401548 420236 401600
rect 421564 401548 421616 401600
rect 433800 401548 433852 401600
rect 341524 401480 341576 401532
rect 347872 401480 347924 401532
rect 353208 401480 353260 401532
rect 443644 401548 443696 401600
rect 451096 401548 451148 401600
rect 472256 401548 472308 401600
rect 449164 401480 449216 401532
rect 334716 401412 334768 401464
rect 370596 401412 370648 401464
rect 323584 401344 323636 401396
rect 440240 401344 440292 401396
rect 447048 401344 447100 401396
rect 482284 401412 482336 401464
rect 324964 401276 325016 401328
rect 443276 401276 443328 401328
rect 446036 401276 446088 401328
rect 472348 401344 472400 401396
rect 472532 401276 472584 401328
rect 342904 401208 342956 401260
rect 346400 401208 346452 401260
rect 353944 401208 353996 401260
rect 360200 401208 360252 401260
rect 362868 401208 362920 401260
rect 480904 401208 480956 401260
rect 327724 401140 327776 401192
rect 354956 401140 355008 401192
rect 478144 401140 478196 401192
rect 322204 401072 322256 401124
rect 350632 401072 350684 401124
rect 356520 401072 356572 401124
rect 476764 401072 476816 401124
rect 343916 401004 343968 401056
rect 474740 401004 474792 401056
rect 316684 400936 316736 400988
rect 455880 400936 455932 400988
rect 472440 400936 472492 400988
rect 316776 400868 316828 400920
rect 456984 400868 457036 400920
rect 478696 400868 478748 400920
rect 530584 400868 530636 400920
rect 344744 400800 344796 400852
rect 409144 400800 409196 400852
rect 410616 400800 410668 400852
rect 427820 400800 427872 400852
rect 431224 400800 431276 400852
rect 436928 400800 436980 400852
rect 453396 400800 453448 400852
rect 472164 400800 472216 400852
rect 349804 400732 349856 400784
rect 363236 400732 363288 400784
rect 363604 400732 363656 400784
rect 418160 400732 418212 400784
rect 331956 400664 332008 400716
rect 364524 400664 364576 400716
rect 372344 400664 372396 400716
rect 382924 400664 382976 400716
rect 408500 400664 408552 400716
rect 417424 400664 417476 400716
rect 430672 400664 430724 400716
rect 359648 400596 359700 400648
rect 370504 400596 370556 400648
rect 382280 400596 382332 400648
rect 395344 400596 395396 400648
rect 414848 400596 414900 400648
rect 399484 400460 399536 400512
rect 411720 400460 411772 400512
rect 413284 400460 413336 400512
rect 424324 400460 424376 400512
rect 407764 400324 407816 400376
rect 421196 400324 421248 400376
rect 472808 400324 472860 400376
rect 476948 400324 477000 400376
rect 364984 400256 365036 400308
rect 366456 400256 366508 400308
rect 393964 400256 394016 400308
rect 402244 400256 402296 400308
rect 472716 400256 472768 400308
rect 474832 400256 474884 400308
rect 365996 400188 366048 400240
rect 367008 400188 367060 400240
rect 369124 400188 369176 400240
rect 369768 400188 369820 400240
rect 371884 400188 371936 400240
rect 372712 400188 372764 400240
rect 374644 400188 374696 400240
rect 375932 400188 375984 400240
rect 378600 400188 378652 400240
rect 379428 400188 379480 400240
rect 388444 400188 388496 400240
rect 392032 400188 392084 400240
rect 396724 400188 396776 400240
rect 398012 400188 398064 400240
rect 403624 400188 403676 400240
rect 404360 400188 404412 400240
rect 410248 400188 410300 400240
rect 411904 400188 411956 400240
rect 413376 400188 413428 400240
rect 414664 400188 414716 400240
rect 422852 400188 422904 400240
rect 423588 400188 423640 400240
rect 432328 400188 432380 400240
rect 433248 400188 433300 400240
rect 435456 400188 435508 400240
rect 436008 400188 436060 400240
rect 458640 400188 458692 400240
rect 459468 400188 459520 400240
rect 472900 400188 472952 400240
rect 473820 400188 473872 400240
rect 475384 400188 475436 400240
rect 476120 400188 476172 400240
rect 479708 400188 479760 400240
rect 480168 400188 480220 400240
rect 462320 400120 462372 400172
rect 463240 400120 463292 400172
rect 467840 400120 467892 400172
rect 468576 400120 468628 400172
rect 320824 397468 320876 397520
rect 337660 397468 337712 397520
rect 322204 396040 322256 396092
rect 337660 396040 337712 396092
rect 482928 395972 482980 396024
rect 536104 395972 536156 396024
rect 329104 394748 329156 394800
rect 337660 394748 337712 394800
rect 321192 394680 321244 394732
rect 337752 394680 337804 394732
rect 330484 393388 330536 393440
rect 337660 393388 337712 393440
rect 323584 393320 323636 393372
rect 337752 393320 337804 393372
rect 331956 392028 332008 392080
rect 337660 392028 337712 392080
rect 325056 391960 325108 392012
rect 337752 391960 337804 392012
rect 482928 391892 482980 391944
rect 529204 391892 529256 391944
rect 334716 390600 334768 390652
rect 337660 390600 337712 390652
rect 324964 390532 325016 390584
rect 337752 390532 337804 390584
rect 328092 389308 328144 389360
rect 337660 389308 337712 389360
rect 327724 389240 327776 389292
rect 337752 389240 337804 389292
rect 322480 389172 322532 389224
rect 337660 389172 337712 389224
rect 316868 389104 316920 389156
rect 337844 389104 337896 389156
rect 318156 389036 318208 389088
rect 337752 389036 337804 389088
rect 328276 387744 328328 387796
rect 337660 387744 337712 387796
rect 329564 387676 329616 387728
rect 337752 387676 337804 387728
rect 325332 386316 325384 386368
rect 337660 386316 337712 386368
rect 482928 386316 482980 386368
rect 533344 386316 533396 386368
rect 330576 386044 330628 386096
rect 337752 386044 337804 386096
rect 320916 384956 320968 385008
rect 337660 384956 337712 385008
rect 322756 384888 322808 384940
rect 337752 384888 337804 384940
rect 322296 383596 322348 383648
rect 337660 383596 337712 383648
rect 334624 383528 334676 383580
rect 337752 383528 337804 383580
rect 331864 382168 331916 382220
rect 336924 382168 336976 382220
rect 482008 382168 482060 382220
rect 538864 382168 538916 382220
rect 330944 382100 330996 382152
rect 337660 382100 337712 382152
rect 323676 380740 323728 380792
rect 337752 380740 337804 380792
rect 319444 380672 319496 380724
rect 336924 380672 336976 380724
rect 329472 379448 329524 379500
rect 337752 379448 337804 379500
rect 319444 378156 319496 378208
rect 337660 378156 337712 378208
rect 482192 378156 482244 378208
rect 580172 378156 580224 378208
rect 328000 378088 328052 378140
rect 337752 378088 337804 378140
rect 482284 378088 482336 378140
rect 580264 378088 580316 378140
rect 318156 376728 318208 376780
rect 337292 376728 337344 376780
rect 318248 376660 318300 376712
rect 337660 376660 337712 376712
rect 330576 375368 330628 375420
rect 337108 375368 337160 375420
rect 318340 375300 318392 375352
rect 337660 375300 337712 375352
rect 318248 374008 318300 374060
rect 337752 374008 337804 374060
rect 322664 373940 322716 373992
rect 337660 373940 337712 373992
rect 326620 372580 326672 372632
rect 337752 372580 337804 372632
rect 482928 372512 482980 372564
rect 537484 372512 537536 372564
rect 318432 371832 318484 371884
rect 337568 371764 337620 371816
rect 318340 371220 318392 371272
rect 336924 371220 336976 371272
rect 321376 371152 321428 371204
rect 337660 371152 337712 371204
rect 318432 369860 318484 369912
rect 337660 369860 337712 369912
rect 322572 369792 322624 369844
rect 337292 369792 337344 369844
rect 333428 368500 333480 368552
rect 337660 368500 337712 368552
rect 318524 368432 318576 368484
rect 337752 368432 337804 368484
rect 329472 367072 329524 367124
rect 337752 367072 337804 367124
rect 335176 365712 335228 365764
rect 337292 365712 337344 365764
rect 332416 365644 332468 365696
rect 337660 365644 337712 365696
rect 328000 364352 328052 364404
rect 337752 364352 337804 364404
rect 482376 364352 482428 364404
rect 580172 364352 580224 364404
rect 335268 364284 335320 364336
rect 337660 364284 337712 364336
rect 322572 362924 322624 362976
rect 337752 362924 337804 362976
rect 328184 362856 328236 362908
rect 337660 362856 337712 362908
rect 322296 361564 322348 361616
rect 337108 361564 337160 361616
rect 325516 361496 325568 361548
rect 336924 361496 336976 361548
rect 329564 360204 329616 360256
rect 337660 360204 337712 360256
rect 319628 359456 319680 359508
rect 337568 359456 337620 359508
rect 320916 358776 320968 358828
rect 337660 358776 337712 358828
rect 335084 358708 335136 358760
rect 336924 358708 336976 358760
rect 325332 357416 325384 357468
rect 337752 357416 337804 357468
rect 319536 357348 319588 357400
rect 337660 357348 337712 357400
rect 332416 354696 332468 354748
rect 337660 354696 337712 354748
rect 330852 354084 330904 354136
rect 337476 354084 337528 354136
rect 334624 353268 334676 353320
rect 337752 353268 337804 353320
rect 329380 353200 329432 353252
rect 337660 353200 337712 353252
rect 331864 351976 331916 352028
rect 337292 351976 337344 352028
rect 323676 351908 323728 351960
rect 336924 351908 336976 351960
rect 326528 351840 326580 351892
rect 337660 351840 337712 351892
rect 330852 350548 330904 350600
rect 337660 350548 337712 350600
rect 332324 350480 332376 350532
rect 337752 350480 337804 350532
rect 328184 349120 328236 349172
rect 337660 349120 337712 349172
rect 324044 349052 324096 349104
rect 337752 349052 337804 349104
rect 334992 347284 335044 347336
rect 337660 347284 337712 347336
rect 325424 347012 325476 347064
rect 336924 347012 336976 347064
rect 325516 346400 325568 346452
rect 337476 346400 337528 346452
rect 330760 346332 330812 346384
rect 337660 346332 337712 346384
rect 334992 345040 335044 345092
rect 337660 345040 337712 345092
rect 318064 344972 318116 345024
rect 337752 344972 337804 345024
rect 324044 343612 324096 343664
rect 337660 343612 337712 343664
rect 333336 343544 333388 343596
rect 337568 343544 337620 343596
rect 329288 343476 329340 343528
rect 337752 343476 337804 343528
rect 336280 342660 336332 342712
rect 336740 342660 336792 342712
rect 322664 342252 322716 342304
rect 337660 342252 337712 342304
rect 333336 339464 333388 339516
rect 337292 339464 337344 339516
rect 332232 339396 332284 339448
rect 337568 339396 337620 339448
rect 332324 338104 332376 338156
rect 337292 338104 337344 338156
rect 326436 338036 326488 338088
rect 337660 338036 337712 338088
rect 326528 336744 326580 336796
rect 337752 336744 337804 336796
rect 321284 336676 321336 336728
rect 337660 336676 337712 336728
rect 330760 335316 330812 335368
rect 337844 335316 337896 335368
rect 323952 335248 324004 335300
rect 337752 335248 337804 335300
rect 321284 333956 321336 334008
rect 337568 333956 337620 334008
rect 323860 333208 323912 333260
rect 337844 333208 337896 333260
rect 329380 332664 329432 332716
rect 337660 332664 337712 332716
rect 323952 332596 324004 332648
rect 337752 332596 337804 332648
rect 332140 332528 332192 332580
rect 337660 332528 337712 332580
rect 160744 331168 160796 331220
rect 161480 331168 161532 331220
rect 176660 331168 176712 331220
rect 322388 331168 322440 331220
rect 337660 331168 337712 331220
rect 334900 331100 334952 331152
rect 337568 331100 337620 331152
rect 335084 329808 335136 329860
rect 337752 329808 337804 329860
rect 325240 329740 325292 329792
rect 337660 329740 337712 329792
rect 332140 328448 332192 328500
rect 337660 328448 337712 328500
rect 322388 327088 322440 327140
rect 337108 327088 337160 327140
rect 330668 327020 330720 327072
rect 337660 327020 337712 327072
rect 331128 325660 331180 325712
rect 337660 325660 337712 325712
rect 321100 325592 321152 325644
rect 337752 325592 337804 325644
rect 482284 325592 482336 325644
rect 580172 325592 580224 325644
rect 318524 324300 318576 324352
rect 337660 324300 337712 324352
rect 329288 322940 329340 322992
rect 337660 322940 337712 322992
rect 156788 322396 156840 322448
rect 337660 322396 337712 322448
rect 278688 322192 278740 322244
rect 336464 322192 336516 322244
rect 179512 321784 179564 321836
rect 223488 321784 223540 321836
rect 179420 321716 179472 321768
rect 226340 321716 226392 321768
rect 51080 321580 51132 321632
rect 62120 321512 62172 321564
rect 62764 321512 62816 321564
rect 179788 321648 179840 321700
rect 228640 321648 228692 321700
rect 229008 321648 229060 321700
rect 204352 321580 204404 321632
rect 231768 321580 231820 321632
rect 337752 321580 337804 321632
rect 180064 321512 180116 321564
rect 327908 321512 327960 321564
rect 336924 321512 336976 321564
rect 71688 321444 71740 321496
rect 337660 321444 337712 321496
rect 63500 321376 63552 321428
rect 63868 321376 63920 321428
rect 178224 321376 178276 321428
rect 179328 321376 179380 321428
rect 219440 321376 219492 321428
rect 220636 321376 220688 321428
rect 246948 321376 247000 321428
rect 326528 321376 326580 321428
rect 179144 321308 179196 321360
rect 220452 321308 220504 321360
rect 253848 321308 253900 321360
rect 334992 321308 335044 321360
rect 178592 321240 178644 321292
rect 203156 321240 203208 321292
rect 241428 321240 241480 321292
rect 323952 321240 324004 321292
rect 117228 321172 117280 321224
rect 329472 321172 329524 321224
rect 89628 321104 89680 321156
rect 332324 321104 332376 321156
rect 86868 321036 86920 321088
rect 330760 321036 330812 321088
rect 84108 320968 84160 321020
rect 329380 320968 329432 321020
rect 77208 320900 77260 320952
rect 331128 320900 331180 320952
rect 81348 320832 81400 320884
rect 336188 320832 336240 320884
rect 60832 320764 60884 320816
rect 178040 320764 178092 320816
rect 179236 320764 179288 320816
rect 211068 320764 211120 320816
rect 143356 320696 143408 320748
rect 232044 320696 232096 320748
rect 143264 320628 143316 320680
rect 233884 320628 233936 320680
rect 66168 320560 66220 320612
rect 179420 320560 179472 320612
rect 179512 320560 179564 320612
rect 215116 320560 215168 320612
rect 19984 320492 20036 320544
rect 63500 320492 63552 320544
rect 179052 320492 179104 320544
rect 216404 320492 216456 320544
rect 19248 320424 19300 320476
rect 62120 320424 62172 320476
rect 178132 320424 178184 320476
rect 178776 320424 178828 320476
rect 216680 320424 216732 320476
rect 179972 320356 180024 320408
rect 218060 320356 218112 320408
rect 60740 320288 60792 320340
rect 178224 320288 178276 320340
rect 179420 320288 179472 320340
rect 179880 320288 179932 320340
rect 202788 320288 202840 320340
rect 56600 320220 56652 320272
rect 19156 320152 19208 320204
rect 65340 320152 65392 320204
rect 66168 320152 66220 320204
rect 18880 320084 18932 320136
rect 44180 320084 44232 320136
rect 51080 320084 51132 320136
rect 79232 320084 79284 320136
rect 157340 320084 157392 320136
rect 19064 320016 19116 320068
rect 50160 320016 50212 320068
rect 51264 320016 51316 320068
rect 77300 320016 77352 320068
rect 176384 320016 176436 320068
rect 18420 319948 18472 320000
rect 59360 319948 59412 320000
rect 78680 319948 78732 320000
rect 177948 320084 178000 320136
rect 180156 320152 180208 320204
rect 204904 320220 204956 320272
rect 208400 320152 208452 320204
rect 19524 319880 19576 319932
rect 75736 319880 75788 319932
rect 179788 320016 179840 320068
rect 200764 320084 200816 320136
rect 204904 320084 204956 320136
rect 224132 320084 224184 320136
rect 334808 320084 334860 320136
rect 337660 320084 337712 320136
rect 236644 320016 236696 320068
rect 178132 319948 178184 320000
rect 19892 319812 19944 319864
rect 66444 319812 66496 319864
rect 74632 319812 74684 319864
rect 179696 319880 179748 319932
rect 178040 319812 178092 319864
rect 211804 319948 211856 320000
rect 229560 319880 229612 319932
rect 271788 319880 271840 319932
rect 322572 319880 322624 319932
rect 18144 319744 18196 319796
rect 73344 319744 73396 319796
rect 179604 319744 179656 319796
rect 19708 319676 19760 319728
rect 68652 319676 68704 319728
rect 70400 319676 70452 319728
rect 176476 319676 176528 319728
rect 176568 319676 176620 319728
rect 18236 319608 18288 319660
rect 72148 319608 72200 319660
rect 178500 319676 178552 319728
rect 211068 319812 211120 319864
rect 221832 319812 221884 319864
rect 222108 319812 222160 319864
rect 277308 319812 277360 319864
rect 333428 319812 333480 319864
rect 210424 319744 210476 319796
rect 269028 319744 269080 319796
rect 329564 319744 329616 319796
rect 179420 319608 179472 319660
rect 180524 319608 180576 319660
rect 207296 319676 207348 319728
rect 208400 319676 208452 319728
rect 222844 319676 222896 319728
rect 274548 319676 274600 319728
rect 335176 319676 335228 319728
rect 17316 319540 17368 319592
rect 71136 319540 71188 319592
rect 179512 319540 179564 319592
rect 231860 319608 231912 319660
rect 264888 319608 264940 319660
rect 332416 319608 332468 319660
rect 18604 319472 18656 319524
rect 52368 319472 52420 319524
rect 178592 319472 178644 319524
rect 213184 319540 213236 319592
rect 233884 319540 233936 319592
rect 303068 319540 303120 319592
rect 231216 319472 231268 319524
rect 231676 319472 231728 319524
rect 232044 319472 232096 319524
rect 302884 319472 302936 319524
rect 19616 319404 19668 319456
rect 53472 319404 53524 319456
rect 179420 319404 179472 319456
rect 179604 319404 179656 319456
rect 233884 319404 233936 319456
rect 256608 319404 256660 319456
rect 336372 319404 336424 319456
rect 18972 319336 19024 319388
rect 59912 319336 59964 319388
rect 178868 319336 178920 319388
rect 18512 319268 18564 319320
rect 50160 319268 50212 319320
rect 178132 319268 178184 319320
rect 178776 319268 178828 319320
rect 40684 319200 40736 319252
rect 176292 319200 176344 319252
rect 176476 319200 176528 319252
rect 179696 319336 179748 319388
rect 234068 319336 234120 319388
rect 179420 319200 179472 319252
rect 179788 319200 179840 319252
rect 235264 319268 235316 319320
rect 238024 319200 238076 319252
rect 42064 319132 42116 319184
rect 178684 319132 178736 319184
rect 201500 319132 201552 319184
rect 202144 319132 202196 319184
rect 202788 319132 202840 319184
rect 225604 319132 225656 319184
rect 20076 319064 20128 319116
rect 36084 319064 36136 319116
rect 196072 319064 196124 319116
rect 211344 319064 211396 319116
rect 37924 318996 37976 319048
rect 197360 318996 197412 319048
rect 18788 318928 18840 318980
rect 39580 318928 39632 318980
rect 198740 318928 198792 318980
rect 231676 318928 231728 318980
rect 316776 318928 316828 318980
rect 36544 318860 36596 318912
rect 195980 318860 196032 318912
rect 224132 318860 224184 318912
rect 316684 318860 316736 318912
rect 18328 318792 18380 318844
rect 45008 318792 45060 318844
rect 204260 318792 204312 318844
rect 228916 318792 228968 318844
rect 337752 318792 337804 318844
rect 176292 318724 176344 318776
rect 176568 318724 176620 318776
rect 281448 318724 281500 318776
rect 326620 318724 326672 318776
rect 259368 318656 259420 318708
rect 330852 318656 330904 318708
rect 251088 318588 251140 318640
rect 322664 318588 322716 318640
rect 326344 318588 326396 318640
rect 337660 318588 337712 318640
rect 249708 318520 249760 318572
rect 333336 318520 333388 318572
rect 222108 318452 222160 318504
rect 323860 318452 323912 318504
rect 207296 318384 207348 318436
rect 330668 318384 330720 318436
rect 179604 318316 179656 318368
rect 179788 318316 179840 318368
rect 203800 318316 203852 318368
rect 334808 318316 334860 318368
rect 159364 318248 159416 318300
rect 336188 318248 336240 318300
rect 99288 318180 99340 318232
rect 328184 318180 328236 318232
rect 93768 318112 93820 318164
rect 324044 318112 324096 318164
rect 91008 318044 91060 318096
rect 336280 318044 336332 318096
rect 68928 317432 68980 317484
rect 336924 317432 336976 317484
rect 156696 317364 156748 317416
rect 337660 317364 337712 317416
rect 226248 316004 226300 316056
rect 337568 316004 337620 316056
rect 329196 315936 329248 315988
rect 337660 315936 337712 315988
rect 238668 315256 238720 315308
rect 335084 315256 335136 315308
rect 223488 314712 223540 314764
rect 337660 314712 337712 314764
rect 66168 314644 66220 314696
rect 337752 314644 337804 314696
rect 156604 314576 156656 314628
rect 337660 314576 337712 314628
rect 64788 313284 64840 313336
rect 337660 313284 337712 313336
rect 325148 313216 325200 313268
rect 337752 313216 337804 313268
rect 482376 313216 482428 313268
rect 580172 313216 580224 313268
rect 219256 312536 219308 312588
rect 327908 312536 327960 312588
rect 222108 311856 222160 311908
rect 337752 311856 337804 311908
rect 178408 311788 178460 311840
rect 337660 311788 337712 311840
rect 62028 310496 62080 310548
rect 337660 310496 337712 310548
rect 332048 310428 332100 310480
rect 337108 310428 337160 310480
rect 219348 309136 219400 309188
rect 337660 309136 337712 309188
rect 173164 309068 173216 309120
rect 337108 309068 337160 309120
rect 59268 307776 59320 307828
rect 337660 307776 337712 307828
rect 170404 307708 170456 307760
rect 337752 307708 337804 307760
rect 216496 306348 216548 306400
rect 337660 306348 337712 306400
rect 321008 306280 321060 306332
rect 337752 306280 337804 306332
rect 56508 304988 56560 305040
rect 337660 304988 337712 305040
rect 169024 304920 169076 304972
rect 337752 304920 337804 304972
rect 213828 303628 213880 303680
rect 337660 303628 337712 303680
rect 333244 303560 333296 303612
rect 336924 303560 336976 303612
rect 53748 302200 53800 302252
rect 337660 302200 337712 302252
rect 166264 302132 166316 302184
rect 337476 302132 337528 302184
rect 16856 301520 16908 301572
rect 17132 301520 17184 301572
rect 177212 301452 177264 301504
rect 211068 300840 211120 300892
rect 337660 300840 337712 300892
rect 327816 300772 327868 300824
rect 337384 300772 337436 300824
rect 52368 299480 52420 299532
rect 337660 299480 337712 299532
rect 162124 299412 162176 299464
rect 337292 299412 337344 299464
rect 16764 298800 16816 298852
rect 17224 298800 17276 298852
rect 177396 298732 177448 298784
rect 209320 298120 209372 298172
rect 337108 298120 337160 298172
rect 200764 298052 200816 298104
rect 336924 298052 336976 298104
rect 202144 297984 202196 298036
rect 337660 297984 337712 298036
rect 178316 296828 178368 296880
rect 197360 296828 197412 296880
rect 178408 296760 178460 296812
rect 198740 296760 198792 296812
rect 48320 296692 48372 296744
rect 337752 296692 337804 296744
rect 197360 296624 197412 296676
rect 337108 296624 337160 296676
rect 198740 296556 198792 296608
rect 337660 296556 337712 296608
rect 238024 295264 238076 295316
rect 337660 295264 337712 295316
rect 239404 294652 239456 294704
rect 316500 294652 316552 294704
rect 220636 294584 220688 294636
rect 321008 294584 321060 294636
rect 178132 293972 178184 294024
rect 204352 293972 204404 294024
rect 316500 293972 316552 294024
rect 336924 293972 336976 294024
rect 3516 293904 3568 293956
rect 327724 293904 327776 293956
rect 235264 293836 235316 293888
rect 337752 293836 337804 293888
rect 236644 293768 236696 293820
rect 337660 293768 337712 293820
rect 303068 293496 303120 293548
rect 327816 293496 327868 293548
rect 266268 293428 266320 293480
rect 325332 293428 325384 293480
rect 204352 293360 204404 293412
rect 325148 293360 325200 293412
rect 213184 293292 213236 293344
rect 336280 293292 336332 293344
rect 114468 293224 114520 293276
rect 328000 293224 328052 293276
rect 234068 292476 234120 292528
rect 337660 292476 337712 292528
rect 233884 292408 233936 292460
rect 337752 292408 337804 292460
rect 262128 292340 262180 292392
rect 323676 292340 323728 292392
rect 244188 292272 244240 292324
rect 321284 292272 321336 292324
rect 237288 292204 237340 292256
rect 322388 292204 322440 292256
rect 220452 292136 220504 292188
rect 322480 292136 322532 292188
rect 216404 292068 216456 292120
rect 332048 292068 332100 292120
rect 96528 292000 96580 292052
rect 325516 292000 325568 292052
rect 78588 291932 78640 291984
rect 332140 291932 332192 291984
rect 19800 291864 19852 291916
rect 20076 291864 20128 291916
rect 73988 291864 74040 291916
rect 329288 291864 329340 291916
rect 206284 291796 206336 291848
rect 329196 291796 329248 291848
rect 284208 291728 284260 291780
rect 330576 291728 330628 291780
rect 195980 291184 196032 291236
rect 196164 291184 196216 291236
rect 106188 291116 106240 291168
rect 336096 291116 336148 291168
rect 102048 291048 102100 291100
rect 331864 291048 331916 291100
rect 104808 290980 104860 291032
rect 334624 290980 334676 291032
rect 140688 290912 140740 290964
rect 157524 290912 157576 290964
rect 316776 290912 316828 290964
rect 337108 290912 337160 290964
rect 111708 290844 111760 290896
rect 322296 290844 322348 290896
rect 118608 290776 118660 290828
rect 318432 290776 318484 290828
rect 121368 290708 121420 290760
rect 318340 290708 318392 290760
rect 122840 290640 122892 290692
rect 318248 290640 318300 290692
rect 126888 290572 126940 290624
rect 318156 290572 318208 290624
rect 139308 290504 139360 290556
rect 157432 290504 157484 290556
rect 157524 290504 157576 290556
rect 299664 290504 299716 290556
rect 317604 290504 317656 290556
rect 318616 290504 318668 290556
rect 151636 290436 151688 290488
rect 160744 290436 160796 290488
rect 157432 290368 157484 290420
rect 299020 290368 299072 290420
rect 310796 290368 310848 290420
rect 317420 290368 317472 290420
rect 318708 290368 318760 290420
rect 232504 290300 232556 290352
rect 337476 290300 337528 290352
rect 234528 290232 234580 290284
rect 318524 290232 318576 290284
rect 286600 290164 286652 290216
rect 319444 290164 319496 290216
rect 108948 290096 109000 290148
rect 320916 290096 320968 290148
rect 178132 289824 178184 289876
rect 204260 289824 204312 289876
rect 204720 289824 204772 289876
rect 229008 289756 229060 289808
rect 337752 289756 337804 289808
rect 229744 289688 229796 289740
rect 337660 289688 337712 289740
rect 299020 289620 299072 289672
rect 317512 289620 317564 289672
rect 327724 289620 327776 289672
rect 302884 289552 302936 289604
rect 318156 289552 318208 289604
rect 222844 289484 222896 289536
rect 317420 289484 317472 289536
rect 215116 289416 215168 289468
rect 322020 289416 322072 289468
rect 16672 289348 16724 289400
rect 70400 289348 70452 289400
rect 217876 289348 217928 289400
rect 324320 289348 324372 289400
rect 17960 289280 18012 289332
rect 74540 289280 74592 289332
rect 204720 289280 204772 289332
rect 331864 289280 331916 289332
rect 17224 289212 17276 289264
rect 77300 289212 77352 289264
rect 177120 289212 177172 289264
rect 337476 289212 337528 289264
rect 17040 289144 17092 289196
rect 336740 289144 336792 289196
rect 17132 289076 17184 289128
rect 78680 289076 78732 289128
rect 318708 289076 318760 289128
rect 338764 289076 338816 289128
rect 180708 289008 180760 289060
rect 195980 289008 196032 289060
rect 178040 288940 178092 288992
rect 196072 288940 196124 288992
rect 177488 288872 177540 288924
rect 337568 288872 337620 288924
rect 177212 288804 177264 288856
rect 337384 288804 337436 288856
rect 177580 288736 177632 288788
rect 177672 288668 177724 288720
rect 338028 288668 338080 288720
rect 177120 288600 177172 288652
rect 177488 288600 177540 288652
rect 177764 288600 177816 288652
rect 337936 288600 337988 288652
rect 177304 288532 177356 288584
rect 337844 288532 337896 288584
rect 177488 288464 177540 288516
rect 177764 288464 177816 288516
rect 177856 288464 177908 288516
rect 336832 288464 336884 288516
rect 160008 288396 160060 288448
rect 320916 288396 320968 288448
rect 225604 288328 225656 288380
rect 336924 288328 336976 288380
rect 226984 288260 227036 288312
rect 337660 288260 337712 288312
rect 227536 288192 227588 288244
rect 337752 288192 337804 288244
rect 211988 287988 212040 288040
rect 337200 287988 337252 288040
rect 211804 287920 211856 287972
rect 337292 287920 337344 287972
rect 36544 287852 36596 287904
rect 209044 287852 209096 287904
rect 334624 287852 334676 287904
rect 19432 287784 19484 287836
rect 37924 287784 37976 287836
rect 210424 287784 210476 287836
rect 337108 287784 337160 287836
rect 19340 287716 19392 287768
rect 40684 287716 40736 287768
rect 195980 287716 196032 287768
rect 337016 287716 337068 287768
rect 18052 287648 18104 287700
rect 42064 287648 42116 287700
rect 196072 287648 196124 287700
rect 337568 287648 337620 287700
rect 336740 287580 336792 287632
rect 337660 287580 337712 287632
rect 16948 287308 17000 287360
rect 150900 287308 150952 287360
rect 151636 287308 151688 287360
rect 180340 287376 180392 287428
rect 180708 287419 180760 287428
rect 180708 287385 180717 287419
rect 180717 287385 180751 287419
rect 180751 287385 180760 287419
rect 180708 287376 180760 287385
rect 318064 287308 318116 287360
rect 157984 287240 158036 287292
rect 177856 287240 177908 287292
rect 322296 287240 322348 287292
rect 337936 287283 337988 287292
rect 337936 287249 337945 287283
rect 337945 287249 337979 287283
rect 337979 287249 337988 287283
rect 337936 287240 337988 287249
rect 338028 287240 338080 287292
rect 337936 287036 337988 287088
rect 338028 287036 338080 287088
rect 19432 286968 19484 287020
rect 316684 286968 316736 287020
rect 317420 286900 317472 286952
rect 19340 286807 19392 286816
rect 19340 286773 19349 286807
rect 19349 286773 19383 286807
rect 19383 286773 19392 286807
rect 19340 286764 19392 286773
rect 336740 286900 336792 286952
rect 337200 286968 337252 287020
rect 336832 286832 336884 286884
rect 337108 286875 337160 286884
rect 337108 286841 337117 286875
rect 337117 286841 337151 286875
rect 337151 286841 337160 286875
rect 337108 286832 337160 286841
rect 337200 286832 337252 286884
rect 338120 286832 338172 286884
rect 337476 286764 337528 286816
rect 337936 286807 337988 286816
rect 337936 286773 337945 286807
rect 337945 286773 337979 286807
rect 337979 286773 337988 286807
rect 337936 286764 337988 286773
rect 337016 285744 337068 285796
rect 337660 285744 337712 285796
rect 336740 285676 336792 285728
rect 337292 285676 337344 285728
rect 322480 285608 322532 285660
rect 337660 285608 337712 285660
rect 323860 285540 323912 285592
rect 337292 285540 337344 285592
rect 336648 285132 336700 285184
rect 337292 285132 337344 285184
rect 337476 284316 337528 284368
rect 337752 284316 337804 284368
rect 321008 284248 321060 284300
rect 337660 284248 337712 284300
rect 327908 284180 327960 284232
rect 337752 284180 337804 284232
rect 178684 283067 178736 283076
rect 178684 283033 178693 283067
rect 178693 283033 178727 283067
rect 178727 283033 178736 283067
rect 178684 283024 178736 283033
rect 178684 282888 178736 282940
rect 324320 282820 324372 282872
rect 337660 282820 337712 282872
rect 332048 282752 332100 282804
rect 337752 282752 337804 282804
rect 337660 282548 337712 282600
rect 337292 282344 337344 282396
rect 337384 282140 337436 282192
rect 322020 281392 322072 281444
rect 337660 281392 337712 281444
rect 334624 278672 334676 278724
rect 337660 278672 337712 278724
rect 330668 278604 330720 278656
rect 337752 278604 337804 278656
rect 337660 278060 337712 278112
rect 338028 278060 338080 278112
rect 337384 277924 337436 277976
rect 338028 277924 338080 277976
rect 337108 277584 337160 277636
rect 337200 277584 337252 277636
rect 19432 277491 19484 277500
rect 19432 277457 19441 277491
rect 19441 277457 19475 277491
rect 19475 277457 19484 277491
rect 19432 277448 19484 277457
rect 337108 277380 337160 277432
rect 337752 277380 337804 277432
rect 19432 277355 19484 277364
rect 19432 277321 19441 277355
rect 19441 277321 19475 277355
rect 19475 277321 19484 277355
rect 19432 277312 19484 277321
rect 331864 277312 331916 277364
rect 337384 277312 337436 277364
rect 329196 277244 329248 277296
rect 337844 277244 337896 277296
rect 325148 275952 325200 276004
rect 337844 275952 337896 276004
rect 334808 275884 334860 275936
rect 337384 275884 337436 275936
rect 322296 274592 322348 274644
rect 337844 274592 337896 274644
rect 482376 273776 482428 273828
rect 485044 273776 485096 273828
rect 318064 273164 318116 273216
rect 337844 273164 337896 273216
rect 482284 273164 482336 273216
rect 580172 273164 580224 273216
rect 319444 271804 319496 271856
rect 337844 271804 337896 271856
rect 323768 271736 323820 271788
rect 337108 271736 337160 271788
rect 320916 270376 320968 270428
rect 337844 270376 337896 270428
rect 178684 267631 178736 267640
rect 178684 267597 178693 267631
rect 178693 267597 178727 267631
rect 178727 267597 178736 267631
rect 178684 267588 178736 267597
rect 481916 264936 481968 264988
rect 483664 264936 483716 264988
rect 327816 262896 327868 262948
rect 336832 262896 336884 262948
rect 337384 262896 337436 262948
rect 318156 262828 318208 262880
rect 337016 262828 337068 262880
rect 337476 262828 337528 262880
rect 319444 262148 319496 262200
rect 319904 262148 319956 262200
rect 319812 261536 319864 261588
rect 337660 261536 337712 261588
rect 319444 261468 319496 261520
rect 337476 261468 337528 261520
rect 319536 260244 319588 260296
rect 337108 260244 337160 260296
rect 319720 260176 319772 260228
rect 337752 260176 337804 260228
rect 319628 260108 319680 260160
rect 337660 260108 337712 260160
rect 318616 259360 318668 259412
rect 337660 259360 337712 259412
rect 482008 259360 482060 259412
rect 580172 259360 580224 259412
rect 327724 259292 327776 259344
rect 336924 259292 336976 259344
rect 338764 258204 338816 258256
rect 340328 258204 340380 258256
rect 19432 258179 19484 258188
rect 19432 258145 19441 258179
rect 19441 258145 19475 258179
rect 19475 258145 19484 258179
rect 19432 258136 19484 258145
rect 178684 258111 178736 258120
rect 178684 258077 178693 258111
rect 178693 258077 178727 258111
rect 178727 258077 178736 258111
rect 178684 258068 178736 258077
rect 19432 258043 19484 258052
rect 19432 258009 19441 258043
rect 19441 258009 19475 258043
rect 19475 258009 19484 258043
rect 19432 258000 19484 258009
rect 179604 258043 179656 258086
rect 179604 258034 179613 258043
rect 179613 258034 179647 258043
rect 179647 258034 179656 258043
rect 336924 258000 336976 258052
rect 339040 258000 339092 258052
rect 178684 257975 178736 257984
rect 178684 257941 178693 257975
rect 178693 257941 178727 257975
rect 178727 257941 178736 257975
rect 178684 257932 178736 257941
rect 179696 257796 179748 257848
rect 336096 256572 336148 256624
rect 345940 256572 345992 256624
rect 347044 256572 347096 256624
rect 365720 256572 365772 256624
rect 327724 256504 327776 256556
rect 361580 256504 361632 256556
rect 331864 256436 331916 256488
rect 367100 256436 367152 256488
rect 367744 256436 367796 256488
rect 369308 256436 369360 256488
rect 374644 256436 374696 256488
rect 390560 256436 390612 256488
rect 334624 256368 334676 256420
rect 379888 256368 379940 256420
rect 320916 256300 320968 256352
rect 350816 256300 350868 256352
rect 352564 256300 352616 256352
rect 408960 256300 409012 256352
rect 475384 256300 475436 256352
rect 477684 256300 477736 256352
rect 340236 256232 340288 256284
rect 397460 256232 397512 256284
rect 318064 256164 318116 256216
rect 405004 256164 405056 256216
rect 322296 256096 322348 256148
rect 415584 256096 415636 256148
rect 436744 256096 436796 256148
rect 473728 256096 473780 256148
rect 323676 256028 323728 256080
rect 455420 256028 455472 256080
rect 324964 255960 325016 256012
rect 463148 255960 463200 256012
rect 465724 255960 465776 256012
rect 475016 255960 475068 256012
rect 340144 255892 340196 255944
rect 344284 255892 344336 255944
rect 339408 255756 339460 255808
rect 340880 255756 340932 255808
rect 341616 255756 341668 255808
rect 370504 255620 370556 255672
rect 373264 255620 373316 255672
rect 345664 255484 345716 255536
rect 348240 255484 348292 255536
rect 338856 255348 338908 255400
rect 346860 255348 346912 255400
rect 179696 253852 179748 253904
rect 179696 253716 179748 253768
rect 336924 253172 336976 253224
rect 337108 253172 337160 253224
rect 459560 253172 459612 253224
rect 460480 253172 460532 253224
rect 179696 244332 179748 244384
rect 177396 244264 177448 244316
rect 177764 244128 177816 244180
rect 179696 244128 179748 244180
rect 179604 243992 179656 244044
rect 19432 238867 19484 238876
rect 19432 238833 19441 238867
rect 19441 238833 19475 238867
rect 19475 238833 19484 238867
rect 19432 238824 19484 238833
rect 19432 238731 19484 238740
rect 19432 238697 19441 238731
rect 19441 238697 19475 238731
rect 19475 238697 19484 238731
rect 19432 238688 19484 238697
rect 179604 234676 179656 234728
rect 179696 234676 179748 234728
rect 179696 234574 179748 234626
rect 482100 233180 482152 233232
rect 579988 233180 580040 233232
rect 179604 225020 179656 225072
rect 179604 224816 179656 224868
rect 319904 223524 319956 223576
rect 336924 223524 336976 223576
rect 158812 220328 158864 220380
rect 160744 220328 160796 220380
rect 19432 219555 19484 219564
rect 19432 219521 19441 219555
rect 19441 219521 19475 219555
rect 19475 219521 19484 219555
rect 19432 219512 19484 219521
rect 19432 219419 19484 219428
rect 19432 219385 19441 219419
rect 19441 219385 19475 219419
rect 19475 219385 19484 219419
rect 19432 219376 19484 219385
rect 482192 219376 482244 219428
rect 580172 219376 580224 219428
rect 158996 218016 159048 218068
rect 160836 218016 160888 218068
rect 179420 215296 179472 215348
rect 179420 215160 179472 215212
rect 157984 211760 158036 211812
rect 177028 211760 177080 211812
rect 179420 210672 179472 210724
rect 178316 210536 178368 210588
rect 179236 210536 179288 210588
rect 179420 210536 179472 210588
rect 179604 210536 179656 210588
rect 178408 210332 178460 210384
rect 179328 210332 179380 210384
rect 179696 210332 179748 210384
rect 19524 209856 19576 209908
rect 19432 209763 19484 209772
rect 19432 209729 19441 209763
rect 19441 209729 19475 209763
rect 19475 209729 19484 209763
rect 19432 209720 19484 209729
rect 19524 209695 19576 209704
rect 19524 209661 19533 209695
rect 19533 209661 19567 209695
rect 19567 209661 19576 209695
rect 19524 209652 19576 209661
rect 19524 209516 19576 209568
rect 19800 209720 19852 209772
rect 19432 209448 19484 209500
rect 19616 209423 19668 209432
rect 19616 209389 19625 209423
rect 19625 209389 19659 209423
rect 19659 209389 19668 209423
rect 19616 209380 19668 209389
rect 19800 209312 19852 209364
rect 178408 205912 178460 205964
rect 178500 205912 178552 205964
rect 178592 205912 178644 205964
rect 178040 205751 178092 205760
rect 178040 205717 178049 205751
rect 178049 205717 178083 205751
rect 178083 205717 178092 205751
rect 178040 205708 178092 205717
rect 179328 205912 179380 205964
rect 179696 205819 179748 205828
rect 179696 205785 179705 205819
rect 179705 205785 179739 205819
rect 179739 205785 179748 205819
rect 179696 205776 179748 205785
rect 178040 205572 178092 205624
rect 178500 205640 178552 205692
rect 178592 205640 178644 205692
rect 178684 205640 178736 205692
rect 179696 205640 179748 205692
rect 159364 204212 159416 204264
rect 160744 204144 160796 204196
rect 177488 204212 177540 204264
rect 160836 204076 160888 204128
rect 177580 204144 177632 204196
rect 17500 204008 17552 204060
rect 177672 204076 177724 204128
rect 17408 203940 17460 203992
rect 20076 203872 20128 203924
rect 159548 203872 159600 203924
rect 318892 204008 318944 204060
rect 317604 203940 317656 203992
rect 17684 203804 17736 203856
rect 317420 203872 317472 203924
rect 318800 203804 318852 203856
rect 3608 203736 3660 203788
rect 331956 203736 332008 203788
rect 30288 203668 30340 203720
rect 370504 203668 370556 203720
rect 27528 203600 27580 203652
rect 367744 203600 367796 203652
rect 106188 203532 106240 203584
rect 458180 203532 458232 203584
rect 17776 203464 17828 203516
rect 317512 203464 317564 203516
rect 17592 203396 17644 203448
rect 177764 203396 177816 203448
rect 179512 203396 179564 203448
rect 16672 203328 16724 203380
rect 69756 203328 69808 203380
rect 159456 203328 159508 203380
rect 176476 203328 176528 203380
rect 17316 203260 17368 203312
rect 71136 203260 71188 203312
rect 177396 203260 177448 203312
rect 180064 203260 180116 203312
rect 231124 203328 231176 203380
rect 229744 203260 229796 203312
rect 18236 203192 18288 203244
rect 72240 203192 72292 203244
rect 178500 203192 178552 203244
rect 232228 203192 232280 203244
rect 19616 203124 19668 203176
rect 75736 203124 75788 203176
rect 179604 203124 179656 203176
rect 233332 203124 233384 203176
rect 18144 203056 18196 203108
rect 73344 203056 73396 203108
rect 178500 203056 178552 203108
rect 179420 203056 179472 203108
rect 234436 203056 234488 203108
rect 17960 202988 18012 203040
rect 74356 202988 74408 203040
rect 179696 202988 179748 203040
rect 235724 202988 235776 203040
rect 17224 202920 17276 202972
rect 76932 202920 76984 202972
rect 177948 202920 178000 202972
rect 238024 202920 238076 202972
rect 17132 202852 17184 202904
rect 78036 202852 78088 202904
rect 176384 202852 176436 202904
rect 237012 202852 237064 202904
rect 17868 202784 17920 202836
rect 157984 202784 158036 202836
rect 3516 202716 3568 202768
rect 334716 202716 334768 202768
rect 119896 202240 119948 202292
rect 436744 202240 436796 202292
rect 23388 202172 23440 202224
rect 347044 202172 347096 202224
rect 113088 202104 113140 202156
rect 465080 202104 465132 202156
rect 17224 201968 17276 202020
rect 17868 201968 17920 202020
rect 19708 201424 19760 201476
rect 67640 201424 67692 201476
rect 79968 201424 80020 201476
rect 157340 201424 157392 201476
rect 179788 201424 179840 201476
rect 224960 201424 225012 201476
rect 238944 201424 238996 201476
rect 316592 201424 316644 201476
rect 19524 201356 19576 201408
rect 37280 201356 37332 201408
rect 179880 201356 179932 201408
rect 223580 201356 223632 201408
rect 302240 201356 302292 201408
rect 303160 201356 303212 201408
rect 336832 201356 336884 201408
rect 19340 201288 19392 201340
rect 36544 201288 36596 201340
rect 179972 201288 180024 201340
rect 222200 201288 222252 201340
rect 302332 201288 302384 201340
rect 303528 201288 303580 201340
rect 337016 201288 337068 201340
rect 19984 201220 20036 201272
rect 63500 201220 63552 201272
rect 180064 201220 180116 201272
rect 195980 201220 196032 201272
rect 19248 201152 19300 201204
rect 62120 201152 62172 201204
rect 179144 201152 179196 201204
rect 219992 201152 220044 201204
rect 18420 201084 18472 201136
rect 59360 201084 59412 201136
rect 179236 201084 179288 201136
rect 219440 201084 219492 201136
rect 18972 201016 19024 201068
rect 59452 201016 59504 201068
rect 179052 201016 179104 201068
rect 215300 201016 215352 201068
rect 18696 200948 18748 201000
rect 55588 200948 55640 201000
rect 178592 200948 178644 201000
rect 211160 200948 211212 201000
rect 19800 200880 19852 200932
rect 52460 200880 52512 200932
rect 143448 200880 143500 200932
rect 302240 200880 302292 200932
rect 18512 200812 18564 200864
rect 51080 200812 51132 200864
rect 178868 200812 178920 200864
rect 211252 200812 211304 200864
rect 18604 200744 18656 200796
rect 51172 200744 51224 200796
rect 143448 200744 143500 200796
rect 302332 200744 302384 200796
rect 19064 200676 19116 200728
rect 49700 200676 49752 200728
rect 178776 200676 178828 200728
rect 209872 200676 209924 200728
rect 18328 200608 18380 200660
rect 44364 200608 44416 200660
rect 178132 200608 178184 200660
rect 204352 200608 204404 200660
rect 18880 200540 18932 200592
rect 44180 200540 44232 200592
rect 178224 200540 178276 200592
rect 204260 200540 204312 200592
rect 18052 200472 18104 200524
rect 41604 200472 41656 200524
rect 176568 200472 176620 200524
rect 200120 200472 200172 200524
rect 20076 200404 20128 200456
rect 40040 200404 40092 200456
rect 178408 200404 178460 200456
rect 201500 200404 201552 200456
rect 18788 200336 18840 200388
rect 38660 200336 38712 200388
rect 178316 200336 178368 200388
rect 198740 200336 198792 200388
rect 19892 200268 19944 200320
rect 66260 200268 66312 200320
rect 178040 200268 178092 200320
rect 197360 200268 197412 200320
rect 19156 200200 19208 200252
rect 64880 200200 64932 200252
rect 178500 200200 178552 200252
rect 196164 200200 196216 200252
rect 201132 200200 201184 200252
rect 201868 200200 201920 200252
rect 19432 200132 19484 200184
rect 35900 200132 35952 200184
rect 178684 200132 178736 200184
rect 220820 200132 220872 200184
rect 482928 193128 482980 193180
rect 580172 193128 580224 193180
rect 3608 188300 3660 188352
rect 330484 188300 330536 188352
rect 482836 179324 482888 179376
rect 580172 179324 580224 179376
rect 482744 153144 482796 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 325056 150356 325108 150408
rect 482652 139340 482704 139392
rect 580172 139340 580224 139392
rect 3516 137232 3568 137284
rect 329104 137232 329156 137284
rect 482560 113092 482612 113144
rect 579804 113092 579856 113144
rect 482468 100648 482520 100700
rect 580172 100648 580224 100700
rect 3240 97928 3292 97980
rect 323584 97928 323636 97980
rect 3608 84804 3660 84856
rect 336004 84804 336056 84856
rect 485044 73108 485096 73160
rect 580172 73108 580224 73160
rect 482376 60664 482428 60716
rect 580172 60664 580224 60716
rect 32404 51824 32456 51876
rect 369860 51824 369912 51876
rect 43444 51756 43496 51808
rect 382280 51756 382332 51808
rect 35164 51688 35216 51740
rect 374000 51688 374052 51740
rect 3424 44820 3476 44872
rect 320824 44820 320876 44872
rect 483664 33056 483716 33108
rect 580172 33056 580224 33108
rect 34428 29860 34480 29912
rect 376760 29860 376812 29912
rect 41328 29792 41380 29844
rect 385040 29792 385092 29844
rect 37188 29724 37240 29776
rect 380900 29724 380952 29776
rect 55128 29656 55180 29708
rect 400220 29656 400272 29708
rect 48228 29588 48280 29640
rect 393320 29588 393372 29640
rect 3516 20612 3568 20664
rect 322204 20612 322256 20664
rect 482284 20612 482336 20664
rect 579988 20612 580040 20664
rect 59268 13268 59320 13320
rect 318064 13268 318116 13320
rect 52368 13200 52420 13252
rect 340236 13200 340288 13252
rect 22744 13132 22796 13184
rect 360200 13132 360252 13184
rect 39304 13064 39356 13116
rect 378140 13064 378192 13116
rect 14464 11704 14516 11756
rect 342260 11704 342312 11756
rect 18604 10480 18656 10532
rect 349160 10480 349212 10532
rect 7564 10412 7616 10464
rect 340880 10412 340932 10464
rect 66168 10344 66220 10396
rect 412640 10344 412692 10396
rect 124128 10276 124180 10328
rect 475384 10276 475436 10328
rect 9956 9188 10008 9240
rect 320916 9188 320968 9240
rect 45468 9120 45520 9172
rect 374644 9120 374696 9172
rect 4068 9052 4120 9104
rect 340144 9052 340196 9104
rect 7656 8984 7708 9036
rect 345664 8984 345716 9036
rect 44272 8916 44324 8968
rect 389180 8916 389232 8968
rect 71504 8236 71556 8288
rect 419540 8236 419592 8288
rect 75000 8168 75052 8220
rect 423680 8168 423732 8220
rect 85672 8100 85724 8152
rect 434720 8100 434772 8152
rect 82084 8032 82136 8084
rect 430580 8032 430632 8084
rect 78588 7964 78640 8016
rect 427820 7964 427872 8016
rect 92756 7896 92808 7948
rect 443000 7896 443052 7948
rect 99840 7828 99892 7880
rect 451280 7828 451332 7880
rect 114008 7760 114060 7812
rect 466460 7760 466512 7812
rect 117596 7692 117648 7744
rect 470600 7692 470652 7744
rect 106924 7624 106976 7676
rect 459652 7624 459704 7676
rect 124680 7556 124732 7608
rect 478880 7556 478932 7608
rect 64328 7488 64380 7540
rect 411260 7488 411312 7540
rect 60832 7420 60884 7472
rect 407120 7420 407172 7472
rect 50160 7352 50212 7404
rect 396080 7352 396132 7404
rect 57244 7284 57296 7336
rect 402980 7284 403032 7336
rect 43076 7216 43128 7268
rect 387800 7216 387852 7268
rect 39580 7148 39632 7200
rect 383660 7148 383712 7200
rect 41880 7080 41932 7132
rect 386420 7080 386472 7132
rect 20628 7012 20680 7064
rect 362960 7012 363012 7064
rect 73804 6808 73856 6860
rect 422300 6808 422352 6860
rect 84476 6740 84528 6792
rect 433340 6740 433392 6792
rect 77392 6672 77444 6724
rect 426440 6672 426492 6724
rect 80888 6604 80940 6656
rect 429292 6604 429344 6656
rect 91560 6536 91612 6588
rect 441620 6536 441672 6588
rect 87972 6468 88024 6520
rect 437480 6468 437532 6520
rect 98644 6400 98696 6452
rect 449900 6400 449952 6452
rect 109316 6332 109368 6384
rect 460940 6332 460992 6384
rect 95148 6264 95200 6316
rect 445760 6264 445812 6316
rect 102232 6196 102284 6248
rect 454040 6196 454092 6248
rect 116400 6128 116452 6180
rect 469220 6128 469272 6180
rect 70308 6060 70360 6112
rect 418160 6060 418212 6112
rect 63224 5992 63276 6044
rect 409880 5992 409932 6044
rect 66720 5924 66772 5976
rect 414020 5924 414072 5976
rect 48964 5856 49016 5908
rect 394700 5856 394752 5908
rect 59636 5788 59688 5840
rect 405740 5788 405792 5840
rect 56048 5720 56100 5772
rect 401600 5720 401652 5772
rect 52552 5652 52604 5704
rect 397552 5652 397604 5704
rect 13544 5584 13596 5636
rect 354680 5584 354732 5636
rect 90364 5448 90416 5500
rect 440240 5448 440292 5500
rect 86868 5380 86920 5432
rect 436100 5380 436152 5432
rect 79692 5312 79744 5364
rect 429200 5312 429252 5364
rect 101036 5244 101088 5296
rect 452660 5244 452712 5296
rect 108120 5176 108172 5228
rect 459560 5176 459612 5228
rect 97448 5108 97500 5160
rect 448520 5108 448572 5160
rect 118792 5040 118844 5092
rect 471980 5040 472032 5092
rect 115204 4972 115256 5024
rect 467840 4972 467892 5024
rect 111616 4904 111668 4956
rect 463700 4904 463752 4956
rect 104532 4836 104584 4888
rect 456800 4836 456852 4888
rect 122288 4768 122340 4820
rect 476120 4768 476172 4820
rect 93952 4700 94004 4752
rect 444380 4700 444432 4752
rect 83280 4632 83332 4684
rect 431960 4632 432012 4684
rect 76196 4564 76248 4616
rect 425060 4564 425112 4616
rect 72608 4496 72660 4548
rect 420920 4496 420972 4548
rect 69112 4428 69164 4480
rect 416780 4428 416832 4480
rect 21824 4360 21876 4412
rect 364340 4360 364392 4412
rect 12348 4292 12400 4344
rect 353300 4292 353352 4344
rect 17040 4224 17092 4276
rect 358820 4224 358872 4276
rect 1676 4088 1728 4140
rect 7564 4088 7616 4140
rect 11152 4088 11204 4140
rect 351920 4088 351972 4140
rect 26516 4020 26568 4072
rect 27528 4020 27580 4072
rect 367192 4020 367244 4072
rect 15936 3952 15988 4004
rect 357440 3952 357492 4004
rect 14740 3884 14792 3936
rect 356060 3884 356112 3936
rect 25320 3816 25372 3868
rect 28908 3816 28960 3868
rect 371240 3816 371292 3868
rect 32404 3748 32456 3800
rect 375380 3748 375432 3800
rect 105728 3680 105780 3732
rect 106188 3680 106240 3732
rect 123484 3680 123536 3732
rect 124128 3680 124180 3732
rect 465724 3680 465776 3732
rect 53748 3612 53800 3664
rect 398840 3612 398892 3664
rect 8760 3544 8812 3596
rect 18604 3544 18656 3596
rect 34796 3544 34848 3596
rect 39304 3544 39356 3596
rect 46664 3544 46716 3596
rect 391940 3544 391992 3596
rect 2872 3476 2924 3528
rect 14464 3476 14516 3528
rect 18236 3476 18288 3528
rect 22744 3476 22796 3528
rect 27712 3476 27764 3528
rect 32312 3476 32364 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 89168 3476 89220 3528
rect 438860 3476 438912 3528
rect 572 3408 624 3460
rect 17224 3408 17276 3460
rect 31300 3408 31352 3460
rect 35164 3408 35216 3460
rect 38384 3408 38436 3460
rect 43444 3408 43496 3460
rect 96252 3408 96304 3460
rect 447140 3408 447192 3460
rect 6460 3340 6512 3392
rect 338856 3340 338908 3392
rect 5264 3272 5316 3324
rect 336096 3272 336148 3324
rect 19432 3068 19484 3120
rect 327724 3204 327776 3256
rect 24216 3136 24268 3188
rect 331864 3136 331916 3188
rect 35992 3068 36044 3120
rect 334624 3068 334676 3120
rect 67916 3000 67968 3052
rect 322296 3000 322348 3052
rect 103336 2932 103388 2984
rect 323676 2932 323728 2984
rect 110512 2864 110564 2916
rect 324964 2864 325016 2916
rect 121092 2796 121144 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 56796 700602 56824 703520
rect 56784 700596 56836 700602
rect 56784 700538 56836 700544
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 121656 702434 121684 703520
rect 121472 702406 121684 702434
rect 105544 700596 105596 700602
rect 105544 700538 105596 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 85486 680096 85542 680105
rect 85486 680031 85542 680040
rect 85500 679046 85528 680031
rect 105556 679946 105584 700538
rect 121472 699802 121500 702406
rect 137848 700602 137876 703520
rect 154132 700670 154160 703520
rect 202800 700738 202828 703520
rect 218992 700806 219020 703520
rect 218980 700800 219032 700806
rect 218980 700742 219032 700748
rect 202788 700732 202840 700738
rect 202788 700674 202840 700680
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 121380 699774 121500 699802
rect 93872 679918 94116 679946
rect 99668 679918 100004 679946
rect 105556 679932 106030 679946
rect 105556 679918 106044 679932
rect 85488 679040 85540 679046
rect 85488 678982 85540 678988
rect 93872 677346 93900 679918
rect 99668 679318 99696 679918
rect 106016 679810 106044 679918
rect 106108 679918 106320 679946
rect 106108 679810 106136 679918
rect 106016 679782 106136 679810
rect 97908 679312 97960 679318
rect 97908 679254 97960 679260
rect 99656 679312 99708 679318
rect 99656 679254 99708 679260
rect 88064 677340 88116 677346
rect 88064 677282 88116 677288
rect 93860 677340 93912 677346
rect 93860 677282 93912 677288
rect 86144 675510 86172 676124
rect 78588 675504 78640 675510
rect 78588 675446 78640 675452
rect 86132 675504 86184 675510
rect 86132 675446 86184 675452
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 78600 632126 78628 675446
rect 82728 672784 82780 672790
rect 82728 672726 82780 672732
rect 78036 632120 78088 632126
rect 78036 632062 78088 632068
rect 78588 632120 78640 632126
rect 78588 632062 78640 632068
rect 78048 629762 78076 632062
rect 82740 629762 82768 672726
rect 88076 634814 88104 677282
rect 90652 676110 90988 676138
rect 96724 676110 96876 676138
rect 90652 672790 90680 676110
rect 96724 672790 96752 676110
rect 90640 672784 90692 672790
rect 90640 672726 90692 672732
rect 92388 672784 92440 672790
rect 92388 672726 92440 672732
rect 96712 672784 96764 672790
rect 96712 672726 96764 672732
rect 87892 634786 88104 634814
rect 87892 629762 87920 634786
rect 77740 629734 78076 629762
rect 82616 629734 82768 629762
rect 87492 629734 87920 629762
rect 92400 629762 92428 672726
rect 97920 634814 97948 679254
rect 97736 634786 97948 634814
rect 102152 676110 102764 676138
rect 97736 629762 97764 634786
rect 92400 629734 92460 629762
rect 97336 629734 97764 629762
rect 102152 629762 102180 676110
rect 106292 654134 106320 679918
rect 108882 676110 108988 676138
rect 106292 654106 106780 654134
rect 106752 629762 106780 654106
rect 108960 632126 108988 676110
rect 111812 654134 111840 679932
rect 121380 679388 121408 699774
rect 251468 699718 251496 703520
rect 267660 700874 267688 703520
rect 283852 700942 283880 703520
rect 316328 702434 316356 703520
rect 316052 702406 316356 702434
rect 283840 700936 283892 700942
rect 283840 700878 283892 700884
rect 267648 700868 267700 700874
rect 267648 700810 267700 700816
rect 250444 699712 250496 699718
rect 250444 699654 250496 699660
rect 251456 699712 251508 699718
rect 251456 699654 251508 699660
rect 250456 680377 250484 699654
rect 316052 682446 316080 702406
rect 332520 701010 332548 703520
rect 332508 701004 332560 701010
rect 332508 700946 332560 700952
rect 348804 700262 348832 703520
rect 348792 700256 348844 700262
rect 348792 700198 348844 700204
rect 397472 700194 397500 703520
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 413664 700126 413692 703520
rect 413652 700120 413704 700126
rect 413652 700062 413704 700068
rect 446140 700058 446168 703520
rect 462228 700528 462280 700534
rect 462228 700470 462280 700476
rect 460940 700392 460992 700398
rect 460940 700334 460992 700340
rect 446128 700052 446180 700058
rect 446128 699994 446180 700000
rect 276296 682440 276348 682446
rect 276296 682382 276348 682388
rect 316040 682440 316092 682446
rect 316040 682382 316092 682388
rect 276308 681766 276336 682382
rect 267188 681760 267240 681766
rect 267188 681702 267240 681708
rect 276296 681760 276348 681766
rect 276296 681702 276348 681708
rect 276756 681760 276808 681766
rect 276756 681702 276808 681708
rect 250442 680368 250498 680377
rect 250442 680303 250498 680312
rect 248432 679918 249458 679946
rect 241426 679552 241482 679561
rect 241426 679487 241482 679496
rect 241440 679318 241468 679487
rect 241428 679312 241480 679318
rect 241428 679254 241480 679260
rect 114756 672586 114784 676124
rect 117700 676110 117990 676138
rect 241454 676110 241560 676138
rect 114744 672580 114796 672586
rect 114744 672522 114796 672528
rect 115848 672580 115900 672586
rect 115848 672522 115900 672528
rect 111812 654106 111932 654134
rect 111904 632738 111932 654106
rect 111892 632732 111944 632738
rect 111892 632674 111944 632680
rect 115860 632126 115888 672522
rect 117700 632738 117728 676110
rect 241532 675510 241560 676110
rect 238668 675504 238720 675510
rect 238668 675446 238720 675452
rect 241520 675504 241572 675510
rect 241520 675446 241572 675452
rect 116584 632732 116636 632738
rect 116584 632674 116636 632680
rect 117688 632732 117740 632738
rect 117688 632674 117740 632680
rect 126428 632732 126480 632738
rect 126428 632674 126480 632680
rect 108948 632120 109000 632126
rect 108948 632062 109000 632068
rect 111800 632120 111852 632126
rect 111800 632062 111852 632068
rect 115848 632120 115900 632126
rect 115848 632062 115900 632068
rect 111812 629762 111840 632062
rect 116596 629762 116624 632674
rect 121552 632120 121604 632126
rect 121552 632062 121604 632068
rect 121564 629762 121592 632062
rect 126440 629762 126468 632674
rect 238680 632126 238708 675446
rect 246316 672110 246344 676124
rect 242808 672104 242860 672110
rect 242808 672046 242860 672052
rect 246304 672104 246356 672110
rect 246304 672046 246356 672052
rect 237932 632120 237984 632126
rect 237932 632062 237984 632068
rect 238668 632120 238720 632126
rect 238668 632062 238720 632068
rect 237944 629762 237972 632062
rect 242820 629762 242848 672046
rect 248432 632330 248460 679918
rect 252204 672110 252232 676124
rect 251180 672104 251232 672110
rect 251180 672046 251232 672052
rect 252192 672104 252244 672110
rect 252192 672046 252244 672052
rect 251192 654134 251220 672046
rect 251192 654106 251956 654134
rect 247684 632324 247736 632330
rect 247684 632266 247736 632272
rect 248420 632324 248472 632330
rect 248420 632266 248472 632272
rect 247696 629762 247724 632266
rect 102152 629734 102212 629762
rect 106752 629734 107180 629762
rect 111812 629734 112056 629762
rect 116596 629734 116932 629762
rect 121564 629734 121900 629762
rect 126440 629734 126776 629762
rect 237636 629734 237972 629762
rect 242512 629734 242848 629762
rect 247388 629734 247724 629762
rect 251928 629762 251956 654106
rect 255332 632126 255360 679932
rect 260852 679918 261142 679946
rect 267200 679932 267228 681702
rect 258244 676110 258580 676138
rect 258552 672110 258580 676110
rect 258540 672104 258592 672110
rect 258540 672046 258592 672052
rect 259368 672104 259420 672110
rect 259368 672046 259420 672052
rect 259380 632126 259408 672046
rect 260852 632194 260880 679918
rect 271880 676320 271932 676326
rect 271880 676262 271932 676268
rect 272892 676320 272944 676326
rect 272944 676268 273286 676274
rect 272892 676262 273286 676268
rect 264224 676110 264652 676138
rect 270112 676110 270448 676138
rect 264624 673454 264652 676110
rect 264624 673426 264928 673454
rect 264900 632874 264928 673426
rect 264888 632868 264940 632874
rect 264888 632810 264940 632816
rect 270420 632806 270448 676110
rect 271892 654134 271920 676262
rect 272904 676246 273286 676262
rect 271892 654106 272012 654134
rect 270408 632800 270460 632806
rect 270408 632742 270460 632748
rect 271984 632738 272012 654106
rect 272064 632868 272116 632874
rect 272064 632810 272116 632816
rect 271972 632732 272024 632738
rect 271972 632674 272024 632680
rect 260840 632188 260892 632194
rect 260840 632130 260892 632136
rect 266728 632188 266780 632194
rect 266728 632130 266780 632136
rect 255320 632120 255372 632126
rect 255320 632062 255372 632068
rect 256884 632120 256936 632126
rect 256884 632062 256936 632068
rect 259368 632120 259420 632126
rect 259368 632062 259420 632068
rect 261760 632120 261812 632126
rect 261760 632062 261812 632068
rect 256896 629762 256924 632062
rect 261772 629762 261800 632062
rect 266740 629762 266768 632130
rect 251928 629734 252356 629762
rect 256896 629734 257232 629762
rect 261772 629734 262108 629762
rect 266740 629734 267076 629762
rect 272076 629626 272104 632810
rect 276768 630034 276796 681702
rect 455328 680400 455380 680406
rect 455328 680342 455380 680348
rect 316684 679312 316736 679318
rect 316684 679254 316736 679260
rect 281540 632800 281592 632806
rect 281540 632742 281592 632748
rect 276768 630006 276842 630034
rect 276814 629748 276842 630006
rect 281552 629762 281580 632742
rect 286324 632732 286376 632738
rect 286324 632674 286376 632680
rect 286336 629762 286364 632674
rect 281552 629734 281796 629762
rect 286336 629734 286672 629762
rect 271952 629598 272104 629626
rect 72792 628312 72844 628318
rect 72792 628254 72844 628260
rect 232872 628312 232924 628318
rect 232872 628254 232924 628260
rect 72700 628244 72752 628250
rect 72700 628186 72752 628192
rect 72608 628108 72660 628114
rect 72608 628050 72660 628056
rect 72620 623529 72648 628050
rect 72606 623520 72662 623529
rect 72606 623455 72662 623464
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3436 422294 3464 606047
rect 3528 576162 3556 619103
rect 72712 602857 72740 628186
rect 72804 615233 72832 628254
rect 130384 628244 130436 628250
rect 130384 628186 130436 628192
rect 232688 628244 232740 628250
rect 232688 628186 232740 628192
rect 73068 628176 73120 628182
rect 73068 628118 73120 628124
rect 72976 627700 73028 627706
rect 72976 627642 73028 627648
rect 72884 627632 72936 627638
rect 72884 627574 72936 627580
rect 72790 615224 72846 615233
rect 72790 615159 72846 615168
rect 72896 611153 72924 627574
rect 72882 611144 72938 611153
rect 72882 611079 72938 611088
rect 72988 606937 73016 627642
rect 73080 619449 73108 628118
rect 74448 628040 74500 628046
rect 74448 627982 74500 627988
rect 74460 627745 74488 627982
rect 74446 627736 74502 627745
rect 74446 627671 74502 627680
rect 129004 627700 129056 627706
rect 129004 627642 129056 627648
rect 73066 619440 73122 619449
rect 73066 619375 73122 619384
rect 129016 607170 129044 627642
rect 129004 607164 129056 607170
rect 129004 607106 129056 607112
rect 72974 606928 73030 606937
rect 72974 606863 73030 606872
rect 130396 603090 130424 628186
rect 130568 628176 130620 628182
rect 130568 628118 130620 628124
rect 130476 627632 130528 627638
rect 130476 627574 130528 627580
rect 130488 611318 130516 627574
rect 130580 619614 130608 628118
rect 133144 628108 133196 628114
rect 133144 628050 133196 628056
rect 133156 623762 133184 628050
rect 133144 623756 133196 623762
rect 133144 623698 133196 623704
rect 130568 619608 130620 619614
rect 130568 619550 130620 619556
rect 232320 619608 232372 619614
rect 232320 619550 232372 619556
rect 232332 619449 232360 619550
rect 232700 619449 232728 628186
rect 232884 628046 232912 628254
rect 289268 628244 289320 628250
rect 289268 628186 289320 628192
rect 233148 628176 233200 628182
rect 233148 628118 233200 628124
rect 232872 628040 232924 628046
rect 232872 627982 232924 627988
rect 233160 627994 233188 628118
rect 235264 628108 235316 628114
rect 235264 628050 235316 628056
rect 235276 628017 235304 628050
rect 235262 628008 235318 628017
rect 232780 627972 232832 627978
rect 232780 627914 232832 627920
rect 232792 623762 232820 627914
rect 232780 623756 232832 623762
rect 232780 623698 232832 623704
rect 232792 623529 232820 623698
rect 232778 623520 232834 623529
rect 232778 623455 232834 623464
rect 232318 619440 232374 619449
rect 232318 619375 232374 619384
rect 232686 619440 232742 619449
rect 232686 619375 232742 619384
rect 232884 615233 232912 627982
rect 233160 627966 233280 627994
rect 233148 627904 233200 627910
rect 233148 627846 233200 627852
rect 233160 627745 233188 627846
rect 233146 627736 233202 627745
rect 233056 627700 233108 627706
rect 233146 627671 233202 627680
rect 233056 627642 233108 627648
rect 232964 627632 233016 627638
rect 232964 627574 233016 627580
rect 232870 615224 232926 615233
rect 232870 615159 232926 615168
rect 232976 611318 233004 627574
rect 130476 611312 130528 611318
rect 130476 611254 130528 611260
rect 232964 611312 233016 611318
rect 232964 611254 233016 611260
rect 232976 611153 233004 611254
rect 232962 611144 233018 611153
rect 232962 611079 233018 611088
rect 232412 607164 232464 607170
rect 232412 607106 232464 607112
rect 232424 606937 232452 607106
rect 233068 606937 233096 627642
rect 233252 627586 233280 627966
rect 235262 627943 235318 627952
rect 289084 627700 289136 627706
rect 289084 627642 289136 627648
rect 233160 627558 233280 627586
rect 232410 606928 232466 606937
rect 232410 606863 232466 606872
rect 233054 606928 233110 606937
rect 233054 606863 233110 606872
rect 233160 603090 233188 627558
rect 289096 606490 289124 627642
rect 289176 627632 289228 627638
rect 289176 627574 289228 627580
rect 289188 610638 289216 627574
rect 289280 618934 289308 628186
rect 290372 628176 290424 628182
rect 290372 628118 290424 628124
rect 290384 625154 290412 628118
rect 290464 628108 290516 628114
rect 290464 628050 290516 628056
rect 290476 627230 290504 628050
rect 313924 628040 313976 628046
rect 313924 627982 313976 627988
rect 290464 627224 290516 627230
rect 290464 627166 290516 627172
rect 290384 625126 290504 625154
rect 289268 618928 289320 618934
rect 289268 618870 289320 618876
rect 289176 610632 289228 610638
rect 289176 610574 289228 610580
rect 289084 606484 289136 606490
rect 289084 606426 289136 606432
rect 130384 603084 130436 603090
rect 130384 603026 130436 603032
rect 233148 603084 233200 603090
rect 233148 603026 233200 603032
rect 233160 602857 233188 603026
rect 72698 602848 72754 602857
rect 72698 602783 72754 602792
rect 233146 602848 233202 602857
rect 233146 602783 233202 602792
rect 290476 602410 290504 625126
rect 313936 614786 313964 627982
rect 313924 614780 313976 614786
rect 313924 614722 313976 614728
rect 290464 602404 290516 602410
rect 290464 602346 290516 602352
rect 72974 598632 73030 598641
rect 72974 598567 73030 598576
rect 231766 598632 231822 598641
rect 231766 598567 231822 598576
rect 72882 594552 72938 594561
rect 72882 594487 72938 594496
rect 72698 586256 72754 586265
rect 72698 586191 72754 586200
rect 71778 577960 71834 577969
rect 71778 577895 71834 577904
rect 71792 576910 71820 577895
rect 17868 576904 17920 576910
rect 17868 576846 17920 576852
rect 71780 576904 71832 576910
rect 71780 576846 71832 576852
rect 72712 576854 72740 586191
rect 72792 582276 72844 582282
rect 72792 582218 72844 582224
rect 72804 577590 72832 582218
rect 72896 577726 72924 594487
rect 72988 582282 73016 598567
rect 73066 590336 73122 590345
rect 73066 590271 73122 590280
rect 72976 582276 73028 582282
rect 72976 582218 73028 582224
rect 73080 582162 73108 590271
rect 72988 582134 73108 582162
rect 72884 577720 72936 577726
rect 72884 577662 72936 577668
rect 72988 577658 73016 582134
rect 73066 582040 73122 582049
rect 73066 581975 73122 581984
rect 72976 577652 73028 577658
rect 72976 577594 73028 577600
rect 72792 577584 72844 577590
rect 72792 577526 72844 577532
rect 73080 577454 73108 581975
rect 231780 577794 231808 598567
rect 233054 594552 233110 594561
rect 233054 594487 233110 594496
rect 232778 590336 232834 590345
rect 232778 590271 232834 590280
rect 231768 577788 231820 577794
rect 231768 577730 231820 577736
rect 231780 577590 231808 577730
rect 232792 577658 232820 590271
rect 232870 586256 232926 586265
rect 232870 586191 232926 586200
rect 232780 577652 232832 577658
rect 232780 577594 232832 577600
rect 231768 577584 231820 577590
rect 75826 577552 75882 577561
rect 231768 577526 231820 577532
rect 75826 577487 75828 577496
rect 75880 577487 75882 577496
rect 75828 577458 75880 577464
rect 73068 577448 73120 577454
rect 73068 577390 73120 577396
rect 3516 576156 3568 576162
rect 3516 576098 3568 576104
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3528 501022 3556 501735
rect 3516 501016 3568 501022
rect 3516 500958 3568 500964
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3528 448594 3556 449511
rect 3516 448588 3568 448594
rect 3516 448530 3568 448536
rect 3436 422266 3556 422294
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3528 409329 3556 422266
rect 3620 409465 3648 514791
rect 3700 409760 3752 409766
rect 3700 409702 3752 409708
rect 3606 409456 3662 409465
rect 3606 409391 3662 409400
rect 3514 409320 3570 409329
rect 3514 409255 3570 409264
rect 3712 406314 3740 409702
rect 3528 406286 3740 406314
rect 3422 405920 3478 405929
rect 3422 405855 3478 405864
rect 3436 345409 3464 405855
rect 3528 397497 3556 406286
rect 3606 406056 3662 406065
rect 3606 405991 3662 406000
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3620 358465 3648 405991
rect 17130 359272 17186 359281
rect 17130 359207 17186 359216
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 17038 332344 17094 332353
rect 17038 332279 17094 332288
rect 17052 330449 17080 332279
rect 17038 330440 17094 330449
rect 17038 330375 17094 330384
rect 3422 321056 3478 321065
rect 3422 320991 3478 321000
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3436 58585 3464 320991
rect 3790 320920 3846 320929
rect 3790 320855 3846 320864
rect 3606 320784 3662 320793
rect 3606 320719 3662 320728
rect 3516 293956 3568 293962
rect 3516 293898 3568 293904
rect 3528 293185 3556 293898
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3514 289096 3570 289105
rect 3514 289031 3570 289040
rect 3528 241097 3556 289031
rect 3620 254153 3648 320719
rect 3804 306241 3832 320855
rect 3790 306232 3846 306241
rect 3790 306167 3846 306176
rect 16856 301572 16908 301578
rect 16856 301514 16908 301520
rect 16764 298852 16816 298858
rect 16764 298794 16816 298800
rect 16672 289400 16724 289406
rect 16672 289342 16724 289348
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3608 203788 3660 203794
rect 3608 203730 3660 203736
rect 3516 202768 3568 202774
rect 3516 202710 3568 202716
rect 3528 201929 3556 202710
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3620 200114 3648 203730
rect 16684 203386 16712 289342
rect 16776 240009 16804 298794
rect 16868 240961 16896 301514
rect 17052 289202 17080 330375
rect 17144 301578 17172 359207
rect 17222 358320 17278 358329
rect 17222 358255 17278 358264
rect 17132 301572 17184 301578
rect 17132 301514 17184 301520
rect 17236 298858 17264 358255
rect 17774 356144 17830 356153
rect 17774 356079 17830 356088
rect 17682 355192 17738 355201
rect 17682 355127 17738 355136
rect 17498 353424 17554 353433
rect 17498 353359 17554 353368
rect 17406 352336 17462 352345
rect 17406 352271 17462 352280
rect 17316 319592 17368 319598
rect 17316 319534 17368 319540
rect 17224 298852 17276 298858
rect 17224 298794 17276 298800
rect 17224 289264 17276 289270
rect 17224 289206 17276 289212
rect 17040 289196 17092 289202
rect 17040 289138 17092 289144
rect 17132 289128 17184 289134
rect 17132 289070 17184 289076
rect 16948 287360 17000 287366
rect 16948 287302 17000 287308
rect 16854 240952 16910 240961
rect 16854 240887 16910 240896
rect 16762 240000 16818 240009
rect 16762 239935 16818 239944
rect 16960 214033 16988 287302
rect 16946 214024 17002 214033
rect 16946 213959 17002 213968
rect 16960 212129 16988 213959
rect 16946 212120 17002 212129
rect 16946 212055 17002 212064
rect 16672 203380 16724 203386
rect 16672 203322 16724 203328
rect 17144 202910 17172 289070
rect 17236 202978 17264 289206
rect 17328 203318 17356 319534
rect 17420 234025 17448 352271
rect 17512 235113 17540 353359
rect 17590 350568 17646 350577
rect 17590 350503 17646 350512
rect 17498 235104 17554 235113
rect 17498 235039 17554 235048
rect 17406 234016 17462 234025
rect 17406 233951 17462 233960
rect 17420 203998 17448 233951
rect 17512 204066 17540 235039
rect 17604 232257 17632 350503
rect 17696 236881 17724 355127
rect 17788 237833 17816 356079
rect 17880 330721 17908 576846
rect 72712 576826 72832 576854
rect 72804 409193 72832 576826
rect 76084 575878 76420 575906
rect 77648 575878 77984 575906
rect 79304 575878 80008 575906
rect 80960 575878 81296 575906
rect 82616 575878 82768 575906
rect 76392 573986 76420 575878
rect 76380 573980 76432 573986
rect 76380 573922 76432 573928
rect 77956 572762 77984 575878
rect 77944 572756 77996 572762
rect 77944 572698 77996 572704
rect 78588 572756 78640 572762
rect 78588 572698 78640 572704
rect 78600 409358 78628 572698
rect 79980 453354 80008 575878
rect 81268 572966 81296 575878
rect 82740 573170 82768 575878
rect 84120 575878 84180 575906
rect 85836 575878 86172 575906
rect 87492 575878 87828 575906
rect 89148 575878 89484 575906
rect 90804 575878 91048 575906
rect 84120 573306 84148 575878
rect 86144 574054 86172 575878
rect 86132 574048 86184 574054
rect 86132 573990 86184 573996
rect 84108 573300 84160 573306
rect 84108 573242 84160 573248
rect 87800 573238 87828 575878
rect 89456 573918 89484 575878
rect 89444 573912 89496 573918
rect 89444 573854 89496 573860
rect 87788 573232 87840 573238
rect 87788 573174 87840 573180
rect 82728 573164 82780 573170
rect 82728 573106 82780 573112
rect 91020 573034 91048 575878
rect 92354 575634 92382 575892
rect 94024 575878 94360 575906
rect 95680 575878 96016 575906
rect 97336 575878 97672 575906
rect 98992 575878 99328 575906
rect 100556 575878 100708 575906
rect 102212 575878 102548 575906
rect 103868 575878 104204 575906
rect 105524 575878 105860 575906
rect 107088 575878 107424 575906
rect 108744 575878 108988 575906
rect 92354 575606 92428 575634
rect 91008 573028 91060 573034
rect 91008 572970 91060 572976
rect 81256 572960 81308 572966
rect 81256 572902 81308 572908
rect 79968 453348 80020 453354
rect 79968 453290 80020 453296
rect 78588 409352 78640 409358
rect 78588 409294 78640 409300
rect 92400 409222 92428 575606
rect 94332 572762 94360 575878
rect 95988 572762 96016 575878
rect 97644 572762 97672 575878
rect 99300 572762 99328 575878
rect 100680 572830 100708 575878
rect 102520 572898 102548 575878
rect 104176 573238 104204 575878
rect 104164 573232 104216 573238
rect 104164 573174 104216 573180
rect 102508 572892 102560 572898
rect 102508 572834 102560 572840
rect 105544 572892 105596 572898
rect 105544 572834 105596 572840
rect 100668 572824 100720 572830
rect 100668 572766 100720 572772
rect 104164 572824 104216 572830
rect 104164 572766 104216 572772
rect 94320 572756 94372 572762
rect 94320 572698 94372 572704
rect 95148 572756 95200 572762
rect 95148 572698 95200 572704
rect 95976 572756 96028 572762
rect 95976 572698 96028 572704
rect 97264 572756 97316 572762
rect 97264 572698 97316 572704
rect 97632 572756 97684 572762
rect 97632 572698 97684 572704
rect 98644 572756 98696 572762
rect 98644 572698 98696 572704
rect 99288 572756 99340 572762
rect 99288 572698 99340 572704
rect 101404 572756 101456 572762
rect 101404 572698 101456 572704
rect 95160 409290 95188 572698
rect 95148 409284 95200 409290
rect 95148 409226 95200 409232
rect 92388 409216 92440 409222
rect 72790 409184 72846 409193
rect 92388 409158 92440 409164
rect 97276 409154 97304 572698
rect 98656 410650 98684 572698
rect 98644 410644 98696 410650
rect 98644 410586 98696 410592
rect 101416 410582 101444 572698
rect 104176 412214 104204 572766
rect 104164 412208 104216 412214
rect 104164 412150 104216 412156
rect 105556 412146 105584 572834
rect 105832 572762 105860 575878
rect 106924 573232 106976 573238
rect 106924 573174 106976 573180
rect 105820 572756 105872 572762
rect 105820 572698 105872 572704
rect 105544 412140 105596 412146
rect 105544 412082 105596 412088
rect 106936 412078 106964 573174
rect 107396 572014 107424 575878
rect 108960 572762 108988 575878
rect 110340 575878 110400 575906
rect 112056 575878 112392 575906
rect 113712 575878 114048 575906
rect 115276 575878 115612 575906
rect 116932 575878 117268 575906
rect 108304 572756 108356 572762
rect 108304 572698 108356 572704
rect 108948 572756 109000 572762
rect 108948 572698 109000 572704
rect 107384 572008 107436 572014
rect 107384 571950 107436 571956
rect 106924 412072 106976 412078
rect 106924 412014 106976 412020
rect 108316 412010 108344 572698
rect 110340 572082 110368 575878
rect 112364 573782 112392 575878
rect 114020 573850 114048 575878
rect 114008 573844 114060 573850
rect 114008 573786 114060 573792
rect 112352 573776 112404 573782
rect 112352 573718 112404 573724
rect 115584 573238 115612 575878
rect 117240 573646 117268 575878
rect 118528 575878 118588 575906
rect 120244 575878 120580 575906
rect 121900 575878 122236 575906
rect 123464 575878 123800 575906
rect 125120 575878 125456 575906
rect 126776 575878 126928 575906
rect 128432 575878 128768 575906
rect 117228 573640 117280 573646
rect 117228 573582 117280 573588
rect 118528 573510 118556 575878
rect 120552 573714 120580 575878
rect 120540 573708 120592 573714
rect 120540 573650 120592 573656
rect 122208 573578 122236 575878
rect 122196 573572 122248 573578
rect 122196 573514 122248 573520
rect 118516 573504 118568 573510
rect 118516 573446 118568 573452
rect 123772 573442 123800 575878
rect 123760 573436 123812 573442
rect 123760 573378 123812 573384
rect 125428 573374 125456 575878
rect 125416 573368 125468 573374
rect 125416 573310 125468 573316
rect 115572 573232 115624 573238
rect 115572 573174 115624 573180
rect 126900 572898 126928 575878
rect 126888 572892 126940 572898
rect 126888 572834 126940 572840
rect 128740 572830 128768 575878
rect 128728 572824 128780 572830
rect 128728 572766 128780 572772
rect 111064 572756 111116 572762
rect 111064 572698 111116 572704
rect 110328 572076 110380 572082
rect 110328 572018 110380 572024
rect 108304 412004 108356 412010
rect 108304 411946 108356 411952
rect 111076 411942 111104 572698
rect 111064 411936 111116 411942
rect 111064 411878 111116 411884
rect 101404 410576 101456 410582
rect 101404 410518 101456 410524
rect 228824 410236 228876 410242
rect 228824 410178 228876 410184
rect 226248 410168 226300 410174
rect 226248 410110 226300 410116
rect 222108 410100 222160 410106
rect 222108 410042 222160 410048
rect 218980 409964 219032 409970
rect 218980 409906 219032 409912
rect 211068 409828 211120 409834
rect 211068 409770 211120 409776
rect 72790 409119 72846 409128
rect 97264 409148 97316 409154
rect 97264 409090 97316 409096
rect 114468 408468 114520 408474
rect 114468 408410 114520 408416
rect 71688 407856 71740 407862
rect 71686 407824 71688 407833
rect 71740 407824 71742 407833
rect 66168 407788 66220 407794
rect 71686 407759 71742 407768
rect 66168 407730 66220 407736
rect 64512 407720 64564 407726
rect 66180 407697 66208 407730
rect 64512 407662 64564 407668
rect 66166 407688 66222 407697
rect 64524 407289 64552 407662
rect 66166 407623 66222 407632
rect 111708 407380 111760 407386
rect 111708 407322 111760 407328
rect 108948 407312 109000 407318
rect 64510 407280 64566 407289
rect 108948 407254 109000 407260
rect 64510 407215 64566 407224
rect 108960 407153 108988 407254
rect 111720 407153 111748 407322
rect 114480 407153 114508 408410
rect 124128 408400 124180 408406
rect 124128 408342 124180 408348
rect 121368 407652 121420 407658
rect 121368 407594 121420 407600
rect 117228 407584 117280 407590
rect 117228 407526 117280 407532
rect 117240 407153 117268 407526
rect 118608 407448 118660 407454
rect 118608 407390 118660 407396
rect 118620 407153 118648 407390
rect 121380 407153 121408 407594
rect 124140 407153 124168 408342
rect 140688 407992 140740 407998
rect 140686 407960 140688 407969
rect 157524 407992 157576 407998
rect 140740 407960 140742 407969
rect 139308 407924 139360 407930
rect 157524 407934 157576 407940
rect 140686 407895 140742 407904
rect 157432 407924 157484 407930
rect 139308 407866 139360 407872
rect 157432 407866 157484 407872
rect 126888 407516 126940 407522
rect 126888 407458 126940 407464
rect 126900 407153 126928 407458
rect 139320 407153 139348 407866
rect 156788 407856 156840 407862
rect 156788 407798 156840 407804
rect 156696 407788 156748 407794
rect 156696 407730 156748 407736
rect 156604 407720 156656 407726
rect 156604 407662 156656 407668
rect 151360 407176 151412 407182
rect 52366 407144 52422 407153
rect 52366 407079 52368 407088
rect 52420 407079 52422 407088
rect 56506 407144 56562 407153
rect 56506 407079 56562 407088
rect 59266 407144 59322 407153
rect 59266 407079 59322 407088
rect 99286 407144 99342 407153
rect 99286 407079 99342 407088
rect 108946 407144 109002 407153
rect 108946 407079 109002 407088
rect 111706 407144 111762 407153
rect 111706 407079 111762 407088
rect 114466 407144 114522 407153
rect 114466 407079 114522 407088
rect 117226 407144 117282 407153
rect 117226 407079 117282 407088
rect 118606 407144 118662 407153
rect 118606 407079 118662 407088
rect 121366 407144 121422 407153
rect 121366 407079 121422 407088
rect 124126 407144 124182 407153
rect 124126 407079 124182 407088
rect 126886 407144 126942 407153
rect 126886 407079 126942 407088
rect 139306 407144 139362 407153
rect 139306 407079 139362 407088
rect 151358 407144 151360 407153
rect 151412 407144 151414 407153
rect 151358 407079 151414 407088
rect 52368 407050 52420 407056
rect 56520 407046 56548 407079
rect 56508 407040 56560 407046
rect 56508 406982 56560 406988
rect 59280 406978 59308 407079
rect 59268 406972 59320 406978
rect 59268 406914 59320 406920
rect 53472 406904 53524 406910
rect 53472 406846 53524 406852
rect 48688 406360 48740 406366
rect 48688 406302 48740 406308
rect 48700 406201 48728 406302
rect 53484 406201 53512 406846
rect 61108 406836 61160 406842
rect 61108 406778 61160 406784
rect 61120 406201 61148 406778
rect 99300 406774 99328 407079
rect 99288 406768 99340 406774
rect 99288 406710 99340 406716
rect 95976 406700 96028 406706
rect 95976 406642 96028 406648
rect 86224 406632 86276 406638
rect 86222 406600 86224 406609
rect 95988 406609 96016 406642
rect 86276 406600 86278 406609
rect 83648 406564 83700 406570
rect 86222 406535 86278 406544
rect 88614 406600 88670 406609
rect 88614 406535 88670 406544
rect 95974 406600 96030 406609
rect 95974 406535 96030 406544
rect 83648 406506 83700 406512
rect 83660 406473 83688 406506
rect 88628 406502 88656 406535
rect 88616 406496 88668 406502
rect 81070 406464 81126 406473
rect 81070 406399 81072 406408
rect 81124 406399 81126 406408
rect 83646 406464 83702 406473
rect 88616 406438 88668 406444
rect 83646 406399 83702 406408
rect 81072 406370 81124 406376
rect 48686 406192 48742 406201
rect 48686 406127 48742 406136
rect 53470 406192 53526 406201
rect 53470 406127 53526 406136
rect 61106 406192 61162 406201
rect 61106 406127 61162 406136
rect 17866 330712 17922 330721
rect 17866 330647 17922 330656
rect 17774 237824 17830 237833
rect 17774 237759 17830 237768
rect 17682 236872 17738 236881
rect 17682 236807 17738 236816
rect 17590 232248 17646 232257
rect 17590 232183 17646 232192
rect 17500 204060 17552 204066
rect 17500 204002 17552 204008
rect 17408 203992 17460 203998
rect 17408 203934 17460 203940
rect 17604 203454 17632 232183
rect 17696 203862 17724 236807
rect 17684 203856 17736 203862
rect 17684 203798 17736 203804
rect 17788 203522 17816 237759
rect 17880 212401 17908 330647
rect 143354 322008 143410 322017
rect 143354 321943 143410 321952
rect 51080 321632 51132 321638
rect 51080 321574 51132 321580
rect 62762 321600 62818 321609
rect 19430 321192 19486 321201
rect 19430 321127 19486 321136
rect 19248 320476 19300 320482
rect 19248 320418 19300 320424
rect 19156 320204 19208 320210
rect 19156 320146 19208 320152
rect 18880 320136 18932 320142
rect 18880 320078 18932 320084
rect 18420 320000 18472 320006
rect 18420 319942 18472 319948
rect 18144 319796 18196 319802
rect 18144 319738 18196 319744
rect 17960 289332 18012 289338
rect 17960 289274 18012 289280
rect 17866 212392 17922 212401
rect 17866 212327 17922 212336
rect 17776 203516 17828 203522
rect 17776 203458 17828 203464
rect 17592 203448 17644 203454
rect 17592 203390 17644 203396
rect 17316 203312 17368 203318
rect 17316 203254 17368 203260
rect 17224 202972 17276 202978
rect 17224 202914 17276 202920
rect 17132 202904 17184 202910
rect 17132 202846 17184 202852
rect 17880 202842 17908 212327
rect 17972 203046 18000 289274
rect 18052 287700 18104 287706
rect 18052 287642 18104 287648
rect 17960 203040 18012 203046
rect 17960 202982 18012 202988
rect 17868 202836 17920 202842
rect 17868 202778 17920 202784
rect 17880 202026 17908 202778
rect 17224 202020 17276 202026
rect 17224 201962 17276 201968
rect 17868 202020 17920 202026
rect 17868 201962 17920 201968
rect 3528 200086 3648 200114
rect 3528 188873 3556 200086
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3608 188352 3660 188358
rect 3608 188294 3660 188300
rect 3516 137284 3568 137290
rect 3516 137226 3568 137232
rect 3528 84697 3556 137226
rect 3620 136785 3648 188294
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 3608 84856 3660 84862
rect 3608 84798 3660 84804
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3620 45529 3648 84798
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 3424 44872 3476 44878
rect 3424 44814 3476 44820
rect 3436 6497 3464 44814
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 4082
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 480 2912 3470
rect 4080 480 4108 9046
rect 7576 4146 7604 10406
rect 9956 9240 10008 9246
rect 9956 9182 10008 9188
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 5264 3324 5316 3330
rect 5264 3266 5316 3272
rect 5276 480 5304 3266
rect 6472 480 6500 3334
rect 7668 480 7696 8978
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 480 8800 3538
rect 9968 480 9996 9182
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 12348 4344 12400 4350
rect 12348 4286 12400 4292
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 480 11192 4082
rect 12360 480 12388 4286
rect 13556 480 13584 5578
rect 14476 3534 14504 11698
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14752 480 14780 3878
rect 15948 480 15976 3946
rect 17052 480 17080 4218
rect 17236 3466 17264 201962
rect 18064 200530 18092 287642
rect 18156 203114 18184 319738
rect 18236 319660 18288 319666
rect 18236 319602 18288 319608
rect 18248 203250 18276 319602
rect 18328 318844 18380 318850
rect 18328 318786 18380 318792
rect 18236 203244 18288 203250
rect 18236 203186 18288 203192
rect 18144 203108 18196 203114
rect 18144 203050 18196 203056
rect 18340 200666 18368 318786
rect 18432 201142 18460 319942
rect 18694 319696 18750 319705
rect 18694 319631 18750 319640
rect 18604 319524 18656 319530
rect 18604 319466 18656 319472
rect 18512 319320 18564 319326
rect 18512 319262 18564 319268
rect 18420 201136 18472 201142
rect 18420 201078 18472 201084
rect 18524 200870 18552 319262
rect 18512 200864 18564 200870
rect 18512 200806 18564 200812
rect 18616 200802 18644 319466
rect 18708 201006 18736 319631
rect 18788 318980 18840 318986
rect 18788 318922 18840 318928
rect 18696 201000 18748 201006
rect 18696 200942 18748 200948
rect 18604 200796 18656 200802
rect 18604 200738 18656 200744
rect 18328 200660 18380 200666
rect 18328 200602 18380 200608
rect 18052 200524 18104 200530
rect 18052 200466 18104 200472
rect 18800 200394 18828 318922
rect 18892 200598 18920 320078
rect 19064 320068 19116 320074
rect 19064 320010 19116 320016
rect 18972 319388 19024 319394
rect 18972 319330 19024 319336
rect 18984 201074 19012 319330
rect 18972 201068 19024 201074
rect 18972 201010 19024 201016
rect 19076 200734 19104 320010
rect 19064 200728 19116 200734
rect 19064 200670 19116 200676
rect 18880 200592 18932 200598
rect 18880 200534 18932 200540
rect 18788 200388 18840 200394
rect 18788 200330 18840 200336
rect 19168 200258 19196 320146
rect 19260 201210 19288 320418
rect 19444 316169 19472 321127
rect 19984 320544 20036 320550
rect 19984 320486 20036 320492
rect 19524 319932 19576 319938
rect 19524 319874 19576 319880
rect 19430 316160 19486 316169
rect 19430 316095 19486 316104
rect 19432 287836 19484 287842
rect 19432 287778 19484 287784
rect 19340 287768 19392 287774
rect 19340 287710 19392 287716
rect 19352 286906 19380 287710
rect 19444 287026 19472 287778
rect 19432 287020 19484 287026
rect 19432 286962 19484 286968
rect 19352 286878 19472 286906
rect 19340 286816 19392 286822
rect 19340 286758 19392 286764
rect 19352 201346 19380 286758
rect 19444 277506 19472 286878
rect 19432 277500 19484 277506
rect 19432 277442 19484 277448
rect 19432 277364 19484 277370
rect 19432 277306 19484 277312
rect 19444 258194 19472 277306
rect 19432 258188 19484 258194
rect 19432 258130 19484 258136
rect 19432 258052 19484 258058
rect 19432 257994 19484 258000
rect 19444 238882 19472 257994
rect 19432 238876 19484 238882
rect 19432 238818 19484 238824
rect 19432 238740 19484 238746
rect 19432 238682 19484 238688
rect 19444 219570 19472 238682
rect 19432 219564 19484 219570
rect 19432 219506 19484 219512
rect 19432 219428 19484 219434
rect 19432 219370 19484 219376
rect 19444 209778 19472 219370
rect 19536 209914 19564 319874
rect 19892 319864 19944 319870
rect 19892 319806 19944 319812
rect 19708 319728 19760 319734
rect 19708 319670 19760 319676
rect 19616 319456 19668 319462
rect 19616 319398 19668 319404
rect 19524 209908 19576 209914
rect 19524 209850 19576 209856
rect 19432 209772 19484 209778
rect 19628 209774 19656 319398
rect 19432 209714 19484 209720
rect 19536 209746 19656 209774
rect 19536 209710 19564 209746
rect 19524 209704 19576 209710
rect 19720 209681 19748 319670
rect 19798 316296 19854 316305
rect 19798 316231 19854 316240
rect 19812 315897 19840 316231
rect 19798 315888 19854 315897
rect 19798 315823 19854 315832
rect 19798 306640 19854 306649
rect 19798 306575 19854 306584
rect 19812 306241 19840 306575
rect 19798 306232 19854 306241
rect 19798 306167 19854 306176
rect 19798 296984 19854 296993
rect 19798 296919 19854 296928
rect 19812 296585 19840 296919
rect 19798 296576 19854 296585
rect 19798 296511 19854 296520
rect 19800 291916 19852 291922
rect 19800 291858 19852 291864
rect 19812 209778 19840 291858
rect 19800 209772 19852 209778
rect 19800 209714 19852 209720
rect 19524 209646 19576 209652
rect 19706 209672 19762 209681
rect 19706 209607 19762 209616
rect 19524 209568 19576 209574
rect 19524 209510 19576 209516
rect 19432 209500 19484 209506
rect 19432 209442 19484 209448
rect 19340 201340 19392 201346
rect 19340 201282 19392 201288
rect 19248 201204 19300 201210
rect 19248 201146 19300 201152
rect 19156 200252 19208 200258
rect 19156 200194 19208 200200
rect 19444 200190 19472 209442
rect 19536 201414 19564 209510
rect 19616 209432 19668 209438
rect 19616 209374 19668 209380
rect 19706 209400 19762 209409
rect 19628 203182 19656 209374
rect 19706 209335 19762 209344
rect 19800 209364 19852 209370
rect 19616 203176 19668 203182
rect 19616 203118 19668 203124
rect 19720 201482 19748 209335
rect 19800 209306 19852 209312
rect 19708 201476 19760 201482
rect 19708 201418 19760 201424
rect 19524 201408 19576 201414
rect 19524 201350 19576 201356
rect 19812 200938 19840 209306
rect 19800 200932 19852 200938
rect 19800 200874 19852 200880
rect 19904 200326 19932 319806
rect 19996 201278 20024 320486
rect 51092 320142 51120 321574
rect 62120 321564 62172 321570
rect 62762 321535 62764 321544
rect 62120 321506 62172 321512
rect 62816 321535 62818 321544
rect 63866 321600 63922 321609
rect 63866 321535 63922 321544
rect 67638 321600 67694 321609
rect 67638 321535 67694 321544
rect 62764 321506 62816 321512
rect 60832 320816 60884 320822
rect 60832 320758 60884 320764
rect 60740 320340 60792 320346
rect 60740 320282 60792 320288
rect 56600 320272 56652 320278
rect 56600 320214 56652 320220
rect 44180 320136 44232 320142
rect 44178 320104 44180 320113
rect 51080 320136 51132 320142
rect 44232 320104 44234 320113
rect 44178 320039 44234 320048
rect 45006 320104 45062 320113
rect 45006 320039 45062 320048
rect 50158 320104 50214 320113
rect 51080 320078 51132 320084
rect 51262 320104 51318 320113
rect 50158 320039 50160 320048
rect 36082 319968 36138 319977
rect 36082 319903 36138 319912
rect 39578 319968 39634 319977
rect 39578 319903 39634 319912
rect 36096 319122 36124 319903
rect 36542 319152 36598 319161
rect 20076 319116 20128 319122
rect 20076 319058 20128 319064
rect 36084 319116 36136 319122
rect 36542 319087 36598 319096
rect 37922 319152 37978 319161
rect 37922 319087 37978 319096
rect 36084 319058 36136 319064
rect 20088 291922 20116 319058
rect 36556 318918 36584 319087
rect 37936 319054 37964 319087
rect 37924 319048 37976 319054
rect 37924 318990 37976 318996
rect 36544 318912 36596 318918
rect 36544 318854 36596 318860
rect 20076 291916 20128 291922
rect 20076 291858 20128 291864
rect 36556 287910 36584 318854
rect 36544 287904 36596 287910
rect 36544 287846 36596 287852
rect 37936 287842 37964 318990
rect 39592 318986 39620 319903
rect 40682 319288 40738 319297
rect 40682 319223 40684 319232
rect 40736 319223 40738 319232
rect 42062 319288 42118 319297
rect 42062 319223 42118 319232
rect 40684 319194 40736 319200
rect 39580 318980 39632 318986
rect 39580 318922 39632 318928
rect 37924 287836 37976 287842
rect 37924 287778 37976 287784
rect 40696 287774 40724 319194
rect 42076 319190 42104 319223
rect 42064 319184 42116 319190
rect 42064 319126 42116 319132
rect 40684 287768 40736 287774
rect 40684 287710 40736 287716
rect 42076 287706 42104 319126
rect 45020 318850 45048 320039
rect 50212 320039 50214 320048
rect 51262 320039 51264 320048
rect 50160 320010 50212 320016
rect 51316 320039 51318 320048
rect 52366 320104 52422 320113
rect 52366 320039 52422 320048
rect 53470 320104 53526 320113
rect 53470 320039 53526 320048
rect 51264 320010 51316 320016
rect 50172 319326 50200 320010
rect 52380 319530 52408 320039
rect 52368 319524 52420 319530
rect 52368 319466 52420 319472
rect 53484 319462 53512 320039
rect 56506 319696 56562 319705
rect 56612 319682 56640 320214
rect 59358 320104 59414 320113
rect 59358 320039 59414 320048
rect 60646 320104 60702 320113
rect 60752 320090 60780 320282
rect 60702 320062 60780 320090
rect 60646 320039 60702 320048
rect 59372 320006 59400 320039
rect 59360 320000 59412 320006
rect 60844 319977 60872 320758
rect 62132 320482 62160 321506
rect 63880 321434 63908 321535
rect 63500 321428 63552 321434
rect 63500 321370 63552 321376
rect 63868 321428 63920 321434
rect 63868 321370 63920 321376
rect 63512 320550 63540 321370
rect 66168 320612 66220 320618
rect 66168 320554 66220 320560
rect 63500 320544 63552 320550
rect 63500 320486 63552 320492
rect 62120 320476 62172 320482
rect 62120 320418 62172 320424
rect 66180 320210 66208 320554
rect 67652 320521 67680 321535
rect 71688 321496 71740 321502
rect 71688 321438 71740 321444
rect 67638 320512 67694 320521
rect 67638 320447 67694 320456
rect 65340 320204 65392 320210
rect 65340 320146 65392 320152
rect 66168 320204 66220 320210
rect 66168 320146 66220 320152
rect 65352 320113 65380 320146
rect 65338 320104 65394 320113
rect 65338 320039 65394 320048
rect 68650 320104 68706 320113
rect 68650 320039 68706 320048
rect 71134 320104 71190 320113
rect 71134 320039 71190 320048
rect 59360 319942 59412 319948
rect 59910 319968 59966 319977
rect 59910 319903 59966 319912
rect 60830 319968 60886 319977
rect 60830 319903 60886 319912
rect 66442 319968 66498 319977
rect 66442 319903 66498 319912
rect 56562 319654 56640 319682
rect 56506 319631 56562 319640
rect 53472 319456 53524 319462
rect 53472 319398 53524 319404
rect 59924 319394 59952 319903
rect 66456 319870 66484 319903
rect 66444 319864 66496 319870
rect 66444 319806 66496 319812
rect 68664 319734 68692 320039
rect 68652 319728 68704 319734
rect 68652 319670 68704 319676
rect 70400 319728 70452 319734
rect 70400 319670 70452 319676
rect 59912 319388 59964 319394
rect 59912 319330 59964 319336
rect 50160 319320 50212 319326
rect 70412 319297 70440 319670
rect 71148 319598 71176 320039
rect 71136 319592 71188 319598
rect 71136 319534 71188 319540
rect 50160 319262 50212 319268
rect 70398 319288 70454 319297
rect 70398 319223 70454 319232
rect 46202 319152 46258 319161
rect 46202 319087 46258 319096
rect 46216 318889 46244 319087
rect 46202 318880 46258 318889
rect 45008 318844 45060 318850
rect 46202 318815 46258 318824
rect 45008 318786 45060 318792
rect 46216 287745 46244 318815
rect 68928 317484 68980 317490
rect 68928 317426 68980 317432
rect 66168 314696 66220 314702
rect 66168 314638 66220 314644
rect 64788 313336 64840 313342
rect 64788 313278 64840 313284
rect 62028 310548 62080 310554
rect 62028 310490 62080 310496
rect 59268 307828 59320 307834
rect 59268 307770 59320 307776
rect 56508 305040 56560 305046
rect 56508 304982 56560 304988
rect 53748 302252 53800 302258
rect 53748 302194 53800 302200
rect 52368 299532 52420 299538
rect 52368 299474 52420 299480
rect 48320 296744 48372 296750
rect 48320 296686 48372 296692
rect 48332 291145 48360 296686
rect 52380 291145 52408 299474
rect 53760 291145 53788 302194
rect 56520 291145 56548 304982
rect 59280 291145 59308 307770
rect 62040 291145 62068 310490
rect 64800 291145 64828 313278
rect 48318 291136 48374 291145
rect 48318 291071 48374 291080
rect 52366 291136 52422 291145
rect 52366 291071 52422 291080
rect 53746 291136 53802 291145
rect 53746 291071 53802 291080
rect 56506 291136 56562 291145
rect 56506 291071 56562 291080
rect 59266 291136 59322 291145
rect 59266 291071 59322 291080
rect 62026 291136 62082 291145
rect 62026 291071 62082 291080
rect 64786 291136 64842 291145
rect 64786 291071 64842 291080
rect 66180 290737 66208 314638
rect 68940 291145 68968 317426
rect 68926 291136 68982 291145
rect 68926 291071 68982 291080
rect 66166 290728 66222 290737
rect 66166 290663 66222 290672
rect 70412 289406 70440 319223
rect 71700 291145 71728 321438
rect 117228 321224 117280 321230
rect 117228 321166 117280 321172
rect 89628 321156 89680 321162
rect 89628 321098 89680 321104
rect 86868 321088 86920 321094
rect 86868 321030 86920 321036
rect 84108 321020 84160 321026
rect 84108 320962 84160 320968
rect 77208 320952 77260 320958
rect 77208 320894 77260 320900
rect 74630 320512 74686 320521
rect 74630 320447 74686 320456
rect 72146 320104 72202 320113
rect 72146 320039 72202 320048
rect 73342 320104 73398 320113
rect 73342 320039 73398 320048
rect 72160 319666 72188 320039
rect 73356 319802 73384 320039
rect 74644 319870 74672 320447
rect 75734 320104 75790 320113
rect 75734 320039 75790 320048
rect 75748 319938 75776 320039
rect 75736 319932 75788 319938
rect 75736 319874 75788 319880
rect 74632 319864 74684 319870
rect 74632 319806 74684 319812
rect 73344 319796 73396 319802
rect 73344 319738 73396 319744
rect 72148 319660 72200 319666
rect 72148 319602 72200 319608
rect 74644 316034 74672 319806
rect 74552 316006 74672 316034
rect 73988 291916 74040 291922
rect 73988 291858 74040 291864
rect 71686 291136 71742 291145
rect 71686 291071 71742 291080
rect 74000 290329 74028 291858
rect 73986 290320 74042 290329
rect 73986 290255 74042 290264
rect 70400 289400 70452 289406
rect 70400 289342 70452 289348
rect 74552 289338 74580 316006
rect 77220 291145 77248 320894
rect 81348 320884 81400 320890
rect 81348 320826 81400 320832
rect 79232 320136 79284 320142
rect 79230 320104 79232 320113
rect 79284 320104 79286 320113
rect 77300 320068 77352 320074
rect 79230 320039 79286 320048
rect 77300 320010 77352 320016
rect 77312 319297 77340 320010
rect 78680 320000 78732 320006
rect 78680 319942 78732 319948
rect 78692 319705 78720 319942
rect 78678 319696 78734 319705
rect 78678 319631 78734 319640
rect 77298 319288 77354 319297
rect 77298 319223 77354 319232
rect 77206 291136 77262 291145
rect 77206 291071 77262 291080
rect 74540 289332 74592 289338
rect 74540 289274 74592 289280
rect 77312 289270 77340 319223
rect 78588 291984 78640 291990
rect 78588 291926 78640 291932
rect 78600 291145 78628 291926
rect 78586 291136 78642 291145
rect 78586 291071 78642 291080
rect 77300 289264 77352 289270
rect 77300 289206 77352 289212
rect 78692 289134 78720 319631
rect 81360 291145 81388 320826
rect 84120 291145 84148 320962
rect 86880 291145 86908 321030
rect 89640 291145 89668 321098
rect 99288 318232 99340 318238
rect 99288 318174 99340 318180
rect 93768 318164 93820 318170
rect 93768 318106 93820 318112
rect 91008 318096 91060 318102
rect 91008 318038 91060 318044
rect 91020 291145 91048 318038
rect 93780 291145 93808 318106
rect 96528 292052 96580 292058
rect 96528 291994 96580 292000
rect 81346 291136 81402 291145
rect 81346 291071 81402 291080
rect 84106 291136 84162 291145
rect 84106 291071 84162 291080
rect 86866 291136 86922 291145
rect 86866 291071 86922 291080
rect 89626 291136 89682 291145
rect 89626 291071 89682 291080
rect 91006 291136 91062 291145
rect 91006 291071 91062 291080
rect 93766 291136 93822 291145
rect 93766 291071 93822 291080
rect 96540 290193 96568 291994
rect 99300 291145 99328 318174
rect 114468 293276 114520 293282
rect 114468 293218 114520 293224
rect 106188 291168 106240 291174
rect 99286 291136 99342 291145
rect 106186 291136 106188 291145
rect 106240 291136 106242 291145
rect 99286 291071 99342 291080
rect 102048 291100 102100 291106
rect 106186 291071 106242 291080
rect 102048 291042 102100 291048
rect 102060 291009 102088 291042
rect 104808 291032 104860 291038
rect 102046 291000 102102 291009
rect 114480 291009 114508 293218
rect 117240 291145 117268 321166
rect 143368 320754 143396 321943
rect 143356 320748 143408 320754
rect 143356 320690 143408 320696
rect 143264 320680 143316 320686
rect 143264 320622 143316 320628
rect 143276 320521 143304 320622
rect 143262 320512 143318 320521
rect 143262 320447 143318 320456
rect 156616 314634 156644 407662
rect 156708 317422 156736 407730
rect 156800 322454 156828 407798
rect 156788 322448 156840 322454
rect 156788 322390 156840 322396
rect 157340 320136 157392 320142
rect 157340 320078 157392 320084
rect 157352 319025 157380 320078
rect 157338 319016 157394 319025
rect 157338 318951 157394 318960
rect 156696 317416 156748 317422
rect 156696 317358 156748 317364
rect 156604 314628 156656 314634
rect 156604 314570 156656 314576
rect 117226 291136 117282 291145
rect 117226 291071 117282 291080
rect 104808 290974 104860 290980
rect 114466 291000 114522 291009
rect 102046 290935 102102 290944
rect 104820 290737 104848 290974
rect 114466 290935 114522 290944
rect 140688 290964 140740 290970
rect 140688 290906 140740 290912
rect 111708 290896 111760 290902
rect 111706 290864 111708 290873
rect 140700 290873 140728 290906
rect 111760 290864 111762 290873
rect 140686 290864 140742 290873
rect 111706 290799 111762 290808
rect 118608 290828 118660 290834
rect 140686 290799 140742 290808
rect 118608 290770 118660 290776
rect 118620 290737 118648 290770
rect 121368 290760 121420 290766
rect 104806 290728 104862 290737
rect 104806 290663 104862 290672
rect 118606 290728 118662 290737
rect 121368 290702 121420 290708
rect 118606 290663 118662 290672
rect 121380 290329 121408 290702
rect 122840 290692 122892 290698
rect 122840 290634 122892 290640
rect 121366 290320 121422 290329
rect 121366 290255 121422 290264
rect 96526 290184 96582 290193
rect 96526 290119 96582 290128
rect 108948 290148 109000 290154
rect 108948 290090 109000 290096
rect 108960 290057 108988 290090
rect 122852 290057 122880 290634
rect 126888 290624 126940 290630
rect 126888 290566 126940 290572
rect 126900 290465 126928 290566
rect 139308 290556 139360 290562
rect 139308 290498 139360 290504
rect 139320 290465 139348 290498
rect 151636 290488 151688 290494
rect 126886 290456 126942 290465
rect 126886 290391 126942 290400
rect 139306 290456 139362 290465
rect 151636 290430 151688 290436
rect 139306 290391 139362 290400
rect 108946 290048 109002 290057
rect 108946 289983 109002 289992
rect 122838 290048 122894 290057
rect 122838 289983 122894 289992
rect 78680 289128 78732 289134
rect 78680 289070 78732 289076
rect 46202 287736 46258 287745
rect 42064 287700 42116 287706
rect 46202 287671 46258 287680
rect 42064 287642 42116 287648
rect 150898 287464 150954 287473
rect 150898 287399 150954 287408
rect 150912 287366 150940 287399
rect 151648 287366 151676 290430
rect 150900 287360 150952 287366
rect 150900 287302 150952 287308
rect 151636 287360 151688 287366
rect 151636 287302 151688 287308
rect 20076 203924 20128 203930
rect 20076 203866 20128 203872
rect 19984 201272 20036 201278
rect 19984 201214 20036 201220
rect 20088 200462 20116 203866
rect 142066 203824 142122 203833
rect 142066 203759 142122 203768
rect 30288 203720 30340 203726
rect 30288 203662 30340 203668
rect 27528 203652 27580 203658
rect 27528 203594 27580 203600
rect 23388 202224 23440 202230
rect 23388 202166 23440 202172
rect 20076 200456 20128 200462
rect 20076 200398 20128 200404
rect 19892 200320 19944 200326
rect 19892 200262 19944 200268
rect 19432 200184 19484 200190
rect 19432 200126 19484 200132
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 3602 18644 10474
rect 20628 7064 20680 7070
rect 20628 7006 20680 7012
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 18248 480 18276 3470
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19444 480 19472 3062
rect 20640 480 20668 7006
rect 21824 4412 21876 4418
rect 21824 4354 21876 4360
rect 21836 480 21864 4354
rect 22756 3534 22784 13126
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 23400 2774 23428 202166
rect 27540 4078 27568 203594
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 25320 3868 25372 3874
rect 25320 3810 25372 3816
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 23032 2746 23428 2774
rect 23032 480 23060 2746
rect 24228 480 24256 3130
rect 25332 480 25360 3810
rect 26528 480 26556 4014
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27724 480 27752 3470
rect 28920 480 28948 3810
rect 30300 2774 30328 203662
rect 106188 203584 106240 203590
rect 69754 203552 69810 203561
rect 69754 203487 69810 203496
rect 71134 203552 71190 203561
rect 71134 203487 71190 203496
rect 72238 203552 72294 203561
rect 72238 203487 72294 203496
rect 73342 203552 73398 203561
rect 73342 203487 73398 203496
rect 74354 203552 74410 203561
rect 74354 203487 74410 203496
rect 75734 203552 75790 203561
rect 75734 203487 75790 203496
rect 78034 203552 78090 203561
rect 106188 203526 106240 203532
rect 78034 203487 78090 203496
rect 69768 203386 69796 203487
rect 69756 203380 69808 203386
rect 69756 203322 69808 203328
rect 71148 203318 71176 203487
rect 71136 203312 71188 203318
rect 71136 203254 71188 203260
rect 72252 203250 72280 203487
rect 72240 203244 72292 203250
rect 72240 203186 72292 203192
rect 73356 203114 73384 203487
rect 73344 203108 73396 203114
rect 73344 203050 73396 203056
rect 74368 203046 74396 203487
rect 75748 203182 75776 203487
rect 75736 203176 75788 203182
rect 75736 203118 75788 203124
rect 74356 203040 74408 203046
rect 74356 202982 74408 202988
rect 76930 203008 76986 203017
rect 76930 202943 76932 202952
rect 76984 202943 76986 202952
rect 76932 202914 76984 202920
rect 78048 202910 78076 203487
rect 78036 202904 78088 202910
rect 78036 202846 78088 202852
rect 41602 202192 41658 202201
rect 41602 202127 41658 202136
rect 37280 201408 37332 201414
rect 35898 201376 35954 201385
rect 35898 201311 35954 201320
rect 36542 201376 36598 201385
rect 36542 201311 36544 201320
rect 35912 200190 35940 201311
rect 36596 201311 36598 201320
rect 37278 201376 37280 201385
rect 37332 201376 37334 201385
rect 37278 201311 37334 201320
rect 38658 201376 38714 201385
rect 38658 201311 38714 201320
rect 40038 201376 40094 201385
rect 40038 201311 40094 201320
rect 36544 201282 36596 201288
rect 38672 200394 38700 201311
rect 40052 200462 40080 201311
rect 41616 200530 41644 202127
rect 67640 201476 67692 201482
rect 67640 201418 67692 201424
rect 79968 201476 80020 201482
rect 79968 201418 80020 201424
rect 67652 201385 67680 201418
rect 79980 201385 80008 201418
rect 44178 201376 44234 201385
rect 44178 201311 44234 201320
rect 44362 201376 44418 201385
rect 44362 201311 44418 201320
rect 63498 201376 63554 201385
rect 63498 201311 63554 201320
rect 67638 201376 67694 201385
rect 67638 201311 67694 201320
rect 79966 201376 80022 201385
rect 79966 201311 80022 201320
rect 44192 200598 44220 201311
rect 44376 200666 44404 201311
rect 63512 201278 63540 201311
rect 63500 201272 63552 201278
rect 51078 201240 51134 201249
rect 51078 201175 51134 201184
rect 52458 201240 52514 201249
rect 52458 201175 52514 201184
rect 55586 201240 55642 201249
rect 55586 201175 55642 201184
rect 59358 201240 59414 201249
rect 59358 201175 59414 201184
rect 62118 201240 62174 201249
rect 63500 201214 63552 201220
rect 62118 201175 62120 201184
rect 51092 200870 51120 201175
rect 52472 200938 52500 201175
rect 55600 201006 55628 201175
rect 59372 201142 59400 201175
rect 62172 201175 62174 201184
rect 62120 201146 62172 201152
rect 59360 201136 59412 201142
rect 59360 201078 59412 201084
rect 59450 201104 59506 201113
rect 59450 201039 59452 201048
rect 59504 201039 59506 201048
rect 59452 201010 59504 201016
rect 55588 201000 55640 201006
rect 55588 200942 55640 200948
rect 52460 200932 52512 200938
rect 52460 200874 52512 200880
rect 51080 200864 51132 200870
rect 49698 200832 49754 200841
rect 51080 200806 51132 200812
rect 51170 200832 51226 200841
rect 49698 200767 49754 200776
rect 51170 200767 51172 200776
rect 49712 200734 49740 200767
rect 51224 200767 51226 200776
rect 51172 200738 51224 200744
rect 49700 200728 49752 200734
rect 49700 200670 49752 200676
rect 62026 200696 62082 200705
rect 44364 200660 44416 200666
rect 62026 200631 62082 200640
rect 44364 200602 44416 200608
rect 44180 200592 44232 200598
rect 44180 200534 44232 200540
rect 41604 200524 41656 200530
rect 41604 200466 41656 200472
rect 40040 200456 40092 200462
rect 40040 200398 40092 200404
rect 38660 200388 38712 200394
rect 38660 200330 38712 200336
rect 35900 200184 35952 200190
rect 35900 200126 35952 200132
rect 32404 51876 32456 51882
rect 32404 51818 32456 51824
rect 32416 6914 32444 51818
rect 43444 51808 43496 51814
rect 43444 51750 43496 51756
rect 35164 51740 35216 51746
rect 35164 51682 35216 51688
rect 34428 29912 34480 29918
rect 34428 29854 34480 29860
rect 32324 6886 32444 6914
rect 32324 3534 32352 6886
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 30116 2746 30328 2774
rect 30116 480 30144 2746
rect 31312 480 31340 3402
rect 32416 480 32444 3742
rect 34440 3534 34468 29854
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 33612 480 33640 3470
rect 34808 480 34836 3538
rect 35176 3466 35204 51682
rect 41328 29844 41380 29850
rect 41328 29786 41380 29792
rect 37188 29776 37240 29782
rect 37188 29718 37240 29724
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 36004 480 36032 3062
rect 37200 480 37228 29718
rect 39304 13116 39356 13122
rect 39304 13058 39356 13064
rect 39316 3602 39344 13058
rect 39580 7200 39632 7206
rect 39580 7142 39632 7148
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38396 480 38424 3402
rect 39592 480 39620 7142
rect 41340 3534 41368 29786
rect 43076 7268 43128 7274
rect 43076 7210 43128 7216
rect 41880 7132 41932 7138
rect 41880 7074 41932 7080
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 40696 480 40724 3470
rect 41892 480 41920 7074
rect 43088 480 43116 7210
rect 43456 3466 43484 51750
rect 55128 29708 55180 29714
rect 55128 29650 55180 29656
rect 48228 29640 48280 29646
rect 48228 29582 48280 29588
rect 45468 9172 45520 9178
rect 45468 9114 45520 9120
rect 44272 8968 44324 8974
rect 44272 8910 44324 8916
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 44284 480 44312 8910
rect 45480 480 45508 9114
rect 48240 6914 48268 29582
rect 52368 13252 52420 13258
rect 52368 13194 52420 13200
rect 50160 7404 50212 7410
rect 50160 7346 50212 7352
rect 47872 6886 48268 6914
rect 46664 3596 46716 3602
rect 46664 3538 46716 3544
rect 46676 480 46704 3538
rect 47872 480 47900 6886
rect 48964 5908 49016 5914
rect 48964 5850 49016 5856
rect 48976 480 49004 5850
rect 50172 480 50200 7346
rect 52380 3534 52408 13194
rect 55140 6914 55168 29650
rect 59268 13320 59320 13326
rect 59268 13262 59320 13268
rect 57244 7336 57296 7342
rect 57244 7278 57296 7284
rect 54956 6886 55168 6914
rect 52552 5704 52604 5710
rect 52552 5646 52604 5652
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 51368 480 51396 3470
rect 52564 480 52592 5646
rect 53748 3664 53800 3670
rect 53748 3606 53800 3612
rect 53760 480 53788 3606
rect 54956 480 54984 6886
rect 56048 5772 56100 5778
rect 56048 5714 56100 5720
rect 56060 480 56088 5714
rect 57256 480 57284 7278
rect 59280 3534 59308 13262
rect 60832 7472 60884 7478
rect 60832 7414 60884 7420
rect 59636 5840 59688 5846
rect 59636 5782 59688 5788
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 58452 480 58480 3470
rect 59648 480 59676 5782
rect 60844 480 60872 7414
rect 62040 480 62068 200631
rect 66258 200424 66314 200433
rect 66258 200359 66314 200368
rect 66272 200326 66300 200359
rect 66260 200320 66312 200326
rect 64878 200288 64934 200297
rect 66260 200262 66312 200268
rect 64878 200223 64880 200232
rect 64932 200223 64934 200232
rect 64880 200194 64932 200200
rect 66168 10396 66220 10402
rect 66168 10338 66220 10344
rect 64328 7540 64380 7546
rect 64328 7482 64380 7488
rect 63224 6044 63276 6050
rect 63224 5986 63276 5992
rect 63236 480 63264 5986
rect 64340 480 64368 7482
rect 66180 3534 66208 10338
rect 71504 8288 71556 8294
rect 71504 8230 71556 8236
rect 70308 6112 70360 6118
rect 70308 6054 70360 6060
rect 66720 5976 66772 5982
rect 66720 5918 66772 5924
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 65536 480 65564 3470
rect 66732 480 66760 5918
rect 69112 4480 69164 4486
rect 69112 4422 69164 4428
rect 67916 3052 67968 3058
rect 67916 2994 67968 3000
rect 67928 480 67956 2994
rect 69124 480 69152 4422
rect 70320 480 70348 6054
rect 71516 480 71544 8230
rect 75000 8220 75052 8226
rect 75000 8162 75052 8168
rect 73804 6860 73856 6866
rect 73804 6802 73856 6808
rect 72608 4548 72660 4554
rect 72608 4490 72660 4496
rect 72620 480 72648 4490
rect 73816 480 73844 6802
rect 75012 480 75040 8162
rect 85672 8152 85724 8158
rect 85672 8094 85724 8100
rect 82084 8084 82136 8090
rect 82084 8026 82136 8032
rect 78588 8016 78640 8022
rect 78588 7958 78640 7964
rect 77392 6724 77444 6730
rect 77392 6666 77444 6672
rect 76196 4616 76248 4622
rect 76196 4558 76248 4564
rect 76208 480 76236 4558
rect 77404 480 77432 6666
rect 78600 480 78628 7958
rect 80888 6656 80940 6662
rect 80888 6598 80940 6604
rect 79692 5364 79744 5370
rect 79692 5306 79744 5312
rect 79704 480 79732 5306
rect 80900 480 80928 6598
rect 82096 480 82124 8026
rect 84476 6792 84528 6798
rect 84476 6734 84528 6740
rect 83280 4684 83332 4690
rect 83280 4626 83332 4632
rect 83292 480 83320 4626
rect 84488 480 84516 6734
rect 85684 480 85712 8094
rect 92756 7948 92808 7954
rect 92756 7890 92808 7896
rect 91560 6588 91612 6594
rect 91560 6530 91612 6536
rect 87972 6520 88024 6526
rect 87972 6462 88024 6468
rect 86868 5432 86920 5438
rect 86868 5374 86920 5380
rect 86880 480 86908 5374
rect 87984 480 88012 6462
rect 90364 5500 90416 5506
rect 90364 5442 90416 5448
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89180 480 89208 3470
rect 90376 480 90404 5442
rect 91572 480 91600 6530
rect 92768 480 92796 7890
rect 99840 7880 99892 7886
rect 99840 7822 99892 7828
rect 98644 6452 98696 6458
rect 98644 6394 98696 6400
rect 95148 6316 95200 6322
rect 95148 6258 95200 6264
rect 93952 4752 94004 4758
rect 93952 4694 94004 4700
rect 93964 480 93992 4694
rect 95160 480 95188 6258
rect 97448 5160 97500 5166
rect 97448 5102 97500 5108
rect 96252 3460 96304 3466
rect 96252 3402 96304 3408
rect 96264 480 96292 3402
rect 97460 480 97488 5102
rect 98656 480 98684 6394
rect 99852 480 99880 7822
rect 102232 6248 102284 6254
rect 102232 6190 102284 6196
rect 101036 5296 101088 5302
rect 101036 5238 101088 5244
rect 101048 480 101076 5238
rect 102244 480 102272 6190
rect 104532 4888 104584 4894
rect 104532 4830 104584 4836
rect 103336 2984 103388 2990
rect 103336 2926 103388 2932
rect 103348 480 103376 2926
rect 104544 480 104572 4830
rect 106200 3738 106228 203526
rect 119896 202292 119948 202298
rect 119896 202234 119948 202240
rect 113088 202156 113140 202162
rect 113088 202098 113140 202104
rect 106924 7676 106976 7682
rect 106924 7618 106976 7624
rect 105728 3732 105780 3738
rect 105728 3674 105780 3680
rect 106188 3732 106240 3738
rect 106188 3674 106240 3680
rect 105740 480 105768 3674
rect 106936 480 106964 7618
rect 113100 6914 113128 202098
rect 114008 7812 114060 7818
rect 114008 7754 114060 7760
rect 112824 6886 113128 6914
rect 109316 6384 109368 6390
rect 109316 6326 109368 6332
rect 108120 5228 108172 5234
rect 108120 5170 108172 5176
rect 108132 480 108160 5170
rect 109328 480 109356 6326
rect 111616 4956 111668 4962
rect 111616 4898 111668 4904
rect 110512 2916 110564 2922
rect 110512 2858 110564 2864
rect 110524 480 110552 2858
rect 111628 480 111656 4898
rect 112824 480 112852 6886
rect 114020 480 114048 7754
rect 117596 7744 117648 7750
rect 117596 7686 117648 7692
rect 116400 6180 116452 6186
rect 116400 6122 116452 6128
rect 115204 5024 115256 5030
rect 115204 4966 115256 4972
rect 115216 480 115244 4966
rect 116412 480 116440 6122
rect 117608 480 117636 7686
rect 118792 5092 118844 5098
rect 118792 5034 118844 5040
rect 118804 480 118832 5034
rect 119908 480 119936 202234
rect 142080 201249 142108 203759
rect 157352 201482 157380 318951
rect 157444 290562 157472 407866
rect 157536 290970 157564 407934
rect 209504 407720 209556 407726
rect 209504 407662 209556 407668
rect 161480 407176 161532 407182
rect 209516 407153 209544 407662
rect 211080 407153 211108 409770
rect 213828 408740 213880 408746
rect 213828 408682 213880 408688
rect 213840 408513 213868 408682
rect 216588 408672 216640 408678
rect 216588 408614 216640 408620
rect 216600 408513 216628 408614
rect 213826 408504 213882 408513
rect 213826 408439 213882 408448
rect 216586 408504 216642 408513
rect 216586 408439 216642 408448
rect 218992 407153 219020 409906
rect 222120 408377 222148 410042
rect 223488 410032 223540 410038
rect 223488 409974 223540 409980
rect 223500 408377 223528 409974
rect 226260 408513 226288 410110
rect 228836 408513 228864 410178
rect 232884 409426 232912 586191
rect 233068 582162 233096 594487
rect 232976 582134 233096 582162
rect 232976 577726 233004 582134
rect 233054 582040 233110 582049
rect 233054 581975 233110 581984
rect 232964 577720 233016 577726
rect 232964 577662 233016 577668
rect 233068 577454 233096 581975
rect 233146 577960 233202 577969
rect 233146 577895 233202 577904
rect 233160 577522 233188 577895
rect 235262 577552 235318 577561
rect 233148 577516 233200 577522
rect 235262 577487 235264 577496
rect 233148 577458 233200 577464
rect 235316 577487 235318 577496
rect 235264 577458 235316 577464
rect 233056 577448 233108 577454
rect 233056 577390 233108 577396
rect 233068 576230 233096 577390
rect 233056 576224 233108 576230
rect 233056 576166 233108 576172
rect 235980 575878 236316 575906
rect 237544 575878 237880 575906
rect 239200 575878 239536 575906
rect 240856 575878 241468 575906
rect 242512 575878 242848 575906
rect 244076 575878 244228 575906
rect 245732 575878 246068 575906
rect 247388 575878 247724 575906
rect 249044 575878 249748 575906
rect 250700 575878 251128 575906
rect 252264 575878 252508 575906
rect 253920 575878 254256 575906
rect 255576 575878 255912 575906
rect 257232 575878 257568 575906
rect 258888 575878 259408 575906
rect 260452 575878 260788 575906
rect 236288 572626 236316 575878
rect 237852 572762 237880 575878
rect 237840 572756 237892 572762
rect 237840 572698 237892 572704
rect 238668 572756 238720 572762
rect 238668 572698 238720 572704
rect 236276 572620 236328 572626
rect 236276 572562 236328 572568
rect 238680 453422 238708 572698
rect 239508 572558 239536 575878
rect 239496 572552 239548 572558
rect 239496 572494 239548 572500
rect 238668 453416 238720 453422
rect 238668 453358 238720 453364
rect 241440 412634 241468 575878
rect 241348 412606 241468 412634
rect 232872 409420 232924 409426
rect 232872 409362 232924 409368
rect 226246 408504 226302 408513
rect 226246 408439 226302 408448
rect 228822 408504 228878 408513
rect 228822 408439 228878 408448
rect 222106 408368 222162 408377
rect 222106 408303 222162 408312
rect 223486 408368 223542 408377
rect 223486 408303 223542 408312
rect 234528 407992 234580 407998
rect 234528 407934 234580 407940
rect 231768 407788 231820 407794
rect 231768 407730 231820 407736
rect 231780 407153 231808 407730
rect 234540 407153 234568 407934
rect 237288 407856 237340 407862
rect 237288 407798 237340 407804
rect 237300 407153 237328 407798
rect 161480 407118 161532 407124
rect 209502 407144 209558 407153
rect 159362 401704 159418 401713
rect 159362 401639 159418 401648
rect 159086 341728 159142 341737
rect 159086 341663 159142 341672
rect 158718 340096 158774 340105
rect 158718 340031 158774 340040
rect 157524 290964 157576 290970
rect 157524 290906 157576 290912
rect 157536 290562 157564 290906
rect 157432 290556 157484 290562
rect 157432 290498 157484 290504
rect 157524 290556 157576 290562
rect 157524 290498 157576 290504
rect 157444 290426 157472 290498
rect 157432 290420 157484 290426
rect 157432 290362 157484 290368
rect 157984 287292 158036 287298
rect 157984 287234 158036 287240
rect 157996 211818 158024 287234
rect 158732 221785 158760 340031
rect 158810 338736 158866 338745
rect 158810 338671 158866 338680
rect 158718 221776 158774 221785
rect 158718 221711 158774 221720
rect 158824 220425 158852 338671
rect 158994 337240 159050 337249
rect 158994 337175 159050 337184
rect 158902 336016 158958 336025
rect 158902 335951 158958 335960
rect 158810 220416 158866 220425
rect 158810 220351 158812 220360
rect 158864 220351 158866 220360
rect 158812 220322 158864 220328
rect 158824 220291 158852 220322
rect 158916 217705 158944 335951
rect 159008 218929 159036 337175
rect 159100 223417 159128 341663
rect 159376 318306 159404 401639
rect 161492 331226 161520 407118
rect 166264 407108 166316 407114
rect 209502 407079 209558 407088
rect 211066 407144 211122 407153
rect 211066 407079 211122 407088
rect 218978 407144 219034 407153
rect 218978 407079 219034 407088
rect 231766 407144 231822 407153
rect 231766 407079 231822 407088
rect 234526 407144 234582 407153
rect 234526 407079 234582 407088
rect 237286 407144 237342 407153
rect 237286 407079 237342 407088
rect 166264 407050 166316 407056
rect 162124 406360 162176 406366
rect 162124 406302 162176 406308
rect 160744 331220 160796 331226
rect 160744 331162 160796 331168
rect 161480 331220 161532 331226
rect 161480 331162 161532 331168
rect 159364 318300 159416 318306
rect 159364 318242 159416 318248
rect 160756 290494 160784 331162
rect 162136 299470 162164 406302
rect 166276 302190 166304 407050
rect 170404 407040 170456 407046
rect 170404 406982 170456 406988
rect 169024 406904 169076 406910
rect 169024 406846 169076 406852
rect 169036 304978 169064 406846
rect 170416 307766 170444 406982
rect 173164 406972 173216 406978
rect 173164 406914 173216 406920
rect 173176 309126 173204 406914
rect 178408 406836 178460 406842
rect 178408 406778 178460 406784
rect 177210 359272 177266 359281
rect 177210 359207 177266 359216
rect 176660 331220 176712 331226
rect 176660 331162 176712 331168
rect 176672 330857 176700 331162
rect 176658 330848 176714 330857
rect 176658 330783 176714 330792
rect 177118 330440 177174 330449
rect 177118 330375 177174 330384
rect 176384 320068 176436 320074
rect 176384 320010 176436 320016
rect 176292 319252 176344 319258
rect 176292 319194 176344 319200
rect 176304 318782 176332 319194
rect 176292 318776 176344 318782
rect 176292 318718 176344 318724
rect 173164 309120 173216 309126
rect 173164 309062 173216 309068
rect 170404 307760 170456 307766
rect 170404 307702 170456 307708
rect 169024 304972 169076 304978
rect 169024 304914 169076 304920
rect 166264 302184 166316 302190
rect 166264 302126 166316 302132
rect 162124 299464 162176 299470
rect 162124 299406 162176 299412
rect 160744 290488 160796 290494
rect 160744 290430 160796 290436
rect 160008 288448 160060 288454
rect 160008 288390 160060 288396
rect 160020 283257 160048 288390
rect 160006 283248 160062 283257
rect 160006 283183 160062 283192
rect 159086 223408 159142 223417
rect 159086 223343 159142 223352
rect 159362 223408 159418 223417
rect 159362 223343 159418 223352
rect 158994 218920 159050 218929
rect 158994 218855 159050 218864
rect 159008 218074 159036 218855
rect 158996 218068 159048 218074
rect 158996 218010 159048 218016
rect 158902 217696 158958 217705
rect 158902 217631 158958 217640
rect 158916 216753 158944 217631
rect 158902 216744 158958 216753
rect 158902 216679 158958 216688
rect 157984 211812 158036 211818
rect 157984 211754 158036 211760
rect 157996 202842 158024 211754
rect 159376 204270 159404 223343
rect 159454 221776 159510 221785
rect 159454 221711 159510 221720
rect 159364 204264 159416 204270
rect 159364 204206 159416 204212
rect 159468 203386 159496 221711
rect 160744 220380 160796 220386
rect 160744 220322 160796 220328
rect 159546 216744 159602 216753
rect 159546 216679 159602 216688
rect 159560 203930 159588 216679
rect 160756 204202 160784 220322
rect 160836 218068 160888 218074
rect 160836 218010 160888 218016
rect 160744 204196 160796 204202
rect 160744 204138 160796 204144
rect 160848 204134 160876 218010
rect 160836 204128 160888 204134
rect 160836 204070 160888 204076
rect 159548 203924 159600 203930
rect 159548 203866 159600 203872
rect 159456 203380 159508 203386
rect 159456 203322 159508 203328
rect 176396 202910 176424 320010
rect 176476 319728 176528 319734
rect 176476 319670 176528 319676
rect 176568 319728 176620 319734
rect 176568 319670 176620 319676
rect 176488 319258 176516 319670
rect 176476 319252 176528 319258
rect 176476 319194 176528 319200
rect 176488 203386 176516 319194
rect 176580 318782 176608 319670
rect 176568 318776 176620 318782
rect 176568 318718 176620 318724
rect 176476 203380 176528 203386
rect 176476 203322 176528 203328
rect 176384 202904 176436 202910
rect 176384 202846 176436 202852
rect 157984 202836 158036 202842
rect 157984 202778 158036 202784
rect 157340 201476 157392 201482
rect 157340 201418 157392 201424
rect 142066 201240 142122 201249
rect 142066 201175 142122 201184
rect 143446 201240 143502 201249
rect 143446 201175 143502 201184
rect 143460 200938 143488 201175
rect 143448 200932 143500 200938
rect 143448 200874 143500 200880
rect 143446 200832 143502 200841
rect 143446 200767 143448 200776
rect 143500 200767 143502 200776
rect 143448 200738 143500 200744
rect 176580 200530 176608 318718
rect 177132 289270 177160 330375
rect 177224 301510 177252 359207
rect 177394 358320 177450 358329
rect 177394 358255 177450 358264
rect 177212 301504 177264 301510
rect 177212 301446 177264 301452
rect 177120 289264 177172 289270
rect 177120 289206 177172 289212
rect 177224 288862 177252 301446
rect 177408 298790 177436 358255
rect 177854 356144 177910 356153
rect 177854 356079 177910 356088
rect 177762 355192 177818 355201
rect 177762 355127 177818 355136
rect 177670 353424 177726 353433
rect 177670 353359 177726 353368
rect 177578 352336 177634 352345
rect 177578 352271 177634 352280
rect 177486 350568 177542 350577
rect 177486 350503 177542 350512
rect 177396 298784 177448 298790
rect 177396 298726 177448 298732
rect 177408 296714 177436 298726
rect 177316 296686 177436 296714
rect 177212 288856 177264 288862
rect 177212 288798 177264 288804
rect 177120 288652 177172 288658
rect 177120 288594 177172 288600
rect 177132 232257 177160 288594
rect 177224 240961 177252 288798
rect 177316 288590 177344 296686
rect 177500 288930 177528 350503
rect 177488 288924 177540 288930
rect 177488 288866 177540 288872
rect 177500 288658 177528 288866
rect 177592 288794 177620 352271
rect 177580 288788 177632 288794
rect 177580 288730 177632 288736
rect 177488 288652 177540 288658
rect 177488 288594 177540 288600
rect 177304 288584 177356 288590
rect 177304 288526 177356 288532
rect 177210 240952 177266 240961
rect 177210 240887 177266 240896
rect 177316 240009 177344 288526
rect 177488 288516 177540 288522
rect 177488 288458 177540 288464
rect 177394 253872 177450 253881
rect 177394 253807 177450 253816
rect 177408 244322 177436 253807
rect 177396 244316 177448 244322
rect 177396 244258 177448 244264
rect 177394 244080 177450 244089
rect 177394 244015 177450 244024
rect 177302 240000 177358 240009
rect 177302 239935 177358 239944
rect 177408 237833 177436 244015
rect 177394 237824 177450 237833
rect 177394 237759 177450 237768
rect 177118 232248 177174 232257
rect 177118 232183 177174 232192
rect 177026 212392 177082 212401
rect 177026 212327 177082 212336
rect 177040 211818 177068 212327
rect 177028 211812 177080 211818
rect 177028 211754 177080 211760
rect 177408 203318 177436 237759
rect 177500 236881 177528 288458
rect 177486 236872 177542 236881
rect 177486 236807 177542 236816
rect 177500 204270 177528 236807
rect 177592 234025 177620 288730
rect 177684 288726 177712 353359
rect 177672 288720 177724 288726
rect 177672 288662 177724 288668
rect 177684 235113 177712 288662
rect 177776 288658 177804 355127
rect 177764 288652 177816 288658
rect 177764 288594 177816 288600
rect 177776 288522 177804 288594
rect 177868 288522 177896 356079
rect 177946 332344 178002 332353
rect 177946 332279 178002 332288
rect 177960 330449 177988 332279
rect 177946 330440 178002 330449
rect 177946 330375 178002 330384
rect 178224 321428 178276 321434
rect 178224 321370 178276 321376
rect 178130 321328 178186 321337
rect 178130 321263 178186 321272
rect 178040 320816 178092 320822
rect 178040 320758 178092 320764
rect 178052 320657 178080 320758
rect 178038 320648 178094 320657
rect 178038 320583 178094 320592
rect 178144 320482 178172 321263
rect 178132 320476 178184 320482
rect 178132 320418 178184 320424
rect 178236 320346 178264 321370
rect 178224 320340 178276 320346
rect 178224 320282 178276 320288
rect 177948 320136 178000 320142
rect 177948 320078 178000 320084
rect 177764 288516 177816 288522
rect 177764 288458 177816 288464
rect 177856 288516 177908 288522
rect 177856 288458 177908 288464
rect 177868 287994 177896 288458
rect 177776 287966 177896 287994
rect 177776 244297 177804 287966
rect 177856 287292 177908 287298
rect 177856 287234 177908 287240
rect 177762 244288 177818 244297
rect 177762 244223 177818 244232
rect 177764 244180 177816 244186
rect 177764 244122 177816 244128
rect 177670 235104 177726 235113
rect 177670 235039 177726 235048
rect 177578 234016 177634 234025
rect 177578 233951 177634 233960
rect 177488 204264 177540 204270
rect 177488 204206 177540 204212
rect 177592 204202 177620 233951
rect 177580 204196 177632 204202
rect 177580 204138 177632 204144
rect 177684 204134 177712 235039
rect 177776 234705 177804 244122
rect 177762 234696 177818 234705
rect 177762 234631 177818 234640
rect 177762 232248 177818 232257
rect 177762 232183 177818 232192
rect 177672 204128 177724 204134
rect 177672 204070 177724 204076
rect 177776 203454 177804 232183
rect 177868 214033 177896 287234
rect 177854 214024 177910 214033
rect 177854 213959 177910 213968
rect 177868 212129 177896 213959
rect 177854 212120 177910 212129
rect 177854 212055 177910 212064
rect 177764 203448 177816 203454
rect 177764 203390 177816 203396
rect 177396 203312 177448 203318
rect 177396 203254 177448 203260
rect 177960 202978 177988 320078
rect 178132 320000 178184 320006
rect 178132 319942 178184 319948
rect 178040 319864 178092 319870
rect 178040 319806 178092 319812
rect 178052 319433 178080 319806
rect 178038 319424 178094 319433
rect 178038 319359 178094 319368
rect 178144 319326 178172 319942
rect 178132 319320 178184 319326
rect 178132 319262 178184 319268
rect 178420 311846 178448 406778
rect 238574 406600 238630 406609
rect 238574 406535 238630 406544
rect 238588 405958 238616 406535
rect 241348 406026 241376 412606
rect 241428 407924 241480 407930
rect 241428 407866 241480 407872
rect 241440 407153 241468 407866
rect 241426 407144 241482 407153
rect 241426 407079 241482 407088
rect 242820 406094 242848 575878
rect 244200 572490 244228 575878
rect 246040 572762 246068 575878
rect 246028 572756 246080 572762
rect 246028 572698 246080 572704
rect 246948 572756 247000 572762
rect 246948 572698 247000 572704
rect 244188 572484 244240 572490
rect 244188 572426 244240 572432
rect 246960 456210 246988 572698
rect 247696 572694 247724 575878
rect 247684 572688 247736 572694
rect 247684 572630 247736 572636
rect 246948 456204 247000 456210
rect 246948 456146 247000 456152
rect 249720 410514 249748 575878
rect 251100 411262 251128 575878
rect 251088 411256 251140 411262
rect 251088 411198 251140 411204
rect 252480 411194 252508 575878
rect 254228 572354 254256 575878
rect 255884 572762 255912 575878
rect 255872 572756 255924 572762
rect 255872 572698 255924 572704
rect 256608 572756 256660 572762
rect 256608 572698 256660 572704
rect 254216 572348 254268 572354
rect 254216 572290 254268 572296
rect 252468 411188 252520 411194
rect 252468 411130 252520 411136
rect 256620 411126 256648 572698
rect 257540 572422 257568 575878
rect 257528 572416 257580 572422
rect 257528 572358 257580 572364
rect 256608 411120 256660 411126
rect 256608 411062 256660 411068
rect 259380 411058 259408 575878
rect 260760 456142 260788 575878
rect 262094 575634 262122 575892
rect 263764 575878 264100 575906
rect 265420 575878 265756 575906
rect 266984 575878 267688 575906
rect 268640 575878 269068 575906
rect 270296 575878 270448 575906
rect 271952 575878 272288 575906
rect 273608 575878 273944 575906
rect 275172 575878 275508 575906
rect 276828 575878 277348 575906
rect 278484 575878 278728 575906
rect 280140 575878 280476 575906
rect 281796 575878 282132 575906
rect 283360 575878 283696 575906
rect 285016 575878 285628 575906
rect 286672 575878 287008 575906
rect 262094 575606 262168 575634
rect 262140 572286 262168 575606
rect 264072 572762 264100 575878
rect 264060 572756 264112 572762
rect 264060 572698 264112 572704
rect 264888 572756 264940 572762
rect 264888 572698 264940 572704
rect 262128 572280 262180 572286
rect 262128 572222 262180 572228
rect 260748 456136 260800 456142
rect 260748 456078 260800 456084
rect 259368 411052 259420 411058
rect 259368 410994 259420 411000
rect 264900 410990 264928 572698
rect 265728 572218 265756 575878
rect 265716 572212 265768 572218
rect 265716 572154 265768 572160
rect 267660 456074 267688 575878
rect 267648 456068 267700 456074
rect 267648 456010 267700 456016
rect 264888 410984 264940 410990
rect 264888 410926 264940 410932
rect 269040 410922 269068 575878
rect 269028 410916 269080 410922
rect 269028 410858 269080 410864
rect 270420 410786 270448 575878
rect 272260 572762 272288 575878
rect 273916 572762 273944 575878
rect 275480 572762 275508 575878
rect 272248 572756 272300 572762
rect 272248 572698 272300 572704
rect 273168 572756 273220 572762
rect 273168 572698 273220 572704
rect 273904 572756 273956 572762
rect 273904 572698 273956 572704
rect 274548 572756 274600 572762
rect 274548 572698 274600 572704
rect 275468 572756 275520 572762
rect 275468 572698 275520 572704
rect 275928 572756 275980 572762
rect 275928 572698 275980 572704
rect 273180 410854 273208 572698
rect 273168 410848 273220 410854
rect 273168 410790 273220 410796
rect 270408 410780 270460 410786
rect 270408 410722 270460 410728
rect 274560 410718 274588 572698
rect 274548 410712 274600 410718
rect 274548 410654 274600 410660
rect 249708 410508 249760 410514
rect 249708 410450 249760 410456
rect 264888 409692 264940 409698
rect 264888 409634 264940 409640
rect 259368 409080 259420 409086
rect 259368 409022 259420 409028
rect 256608 409012 256660 409018
rect 256608 408954 256660 408960
rect 253848 408876 253900 408882
rect 253848 408818 253900 408824
rect 251088 408808 251140 408814
rect 251088 408750 251140 408756
rect 251100 408513 251128 408750
rect 253860 408513 253888 408818
rect 251086 408504 251142 408513
rect 251086 408439 251142 408448
rect 253846 408504 253902 408513
rect 253846 408439 253902 408448
rect 249708 408128 249760 408134
rect 249708 408070 249760 408076
rect 246948 408060 247000 408066
rect 246948 408002 247000 408008
rect 246960 407153 246988 408002
rect 249720 407153 249748 408070
rect 256620 407153 256648 408954
rect 259380 408513 259408 409022
rect 264900 408513 264928 409634
rect 274548 409556 274600 409562
rect 274548 409498 274600 409504
rect 271788 409488 271840 409494
rect 271788 409430 271840 409436
rect 266268 408944 266320 408950
rect 266268 408886 266320 408892
rect 266280 408513 266308 408886
rect 259366 408504 259422 408513
rect 259366 408439 259422 408448
rect 264886 408504 264942 408513
rect 264886 408439 264942 408448
rect 266266 408504 266322 408513
rect 266266 408439 266322 408448
rect 271800 408377 271828 409430
rect 274560 408513 274588 409498
rect 274546 408504 274602 408513
rect 274546 408439 274602 408448
rect 271786 408368 271842 408377
rect 271786 408303 271842 408312
rect 269028 408264 269080 408270
rect 269028 408206 269080 408212
rect 262128 408196 262180 408202
rect 262128 408138 262180 408144
rect 262140 407153 262168 408138
rect 269040 408105 269068 408206
rect 269026 408096 269082 408105
rect 269026 408031 269082 408040
rect 246946 407144 247002 407153
rect 246946 407079 247002 407088
rect 249706 407144 249762 407153
rect 249706 407079 249762 407088
rect 256606 407144 256662 407153
rect 256606 407079 256662 407088
rect 262126 407144 262182 407153
rect 262126 407079 262182 407088
rect 243726 406600 243782 406609
rect 243726 406535 243782 406544
rect 242808 406088 242860 406094
rect 242808 406030 242860 406036
rect 241336 406020 241388 406026
rect 241336 405962 241388 405968
rect 238576 405952 238628 405958
rect 238576 405894 238628 405900
rect 243740 405890 243768 406535
rect 275940 406162 275968 572698
rect 276848 408536 276900 408542
rect 276848 408478 276900 408484
rect 276860 407153 276888 408478
rect 276846 407144 276902 407153
rect 276846 407079 276902 407088
rect 277320 406230 277348 575878
rect 278700 412634 278728 575878
rect 280448 572762 280476 575878
rect 282104 572762 282132 575878
rect 283668 572762 283696 575878
rect 280436 572756 280488 572762
rect 280436 572698 280488 572704
rect 281448 572756 281500 572762
rect 281448 572698 281500 572704
rect 282092 572756 282144 572762
rect 282092 572698 282144 572704
rect 282828 572756 282880 572762
rect 282828 572698 282880 572704
rect 283656 572756 283708 572762
rect 283656 572698 283708 572704
rect 284208 572756 284260 572762
rect 284208 572698 284260 572704
rect 278608 412606 278728 412634
rect 278608 406298 278636 412606
rect 278688 409624 278740 409630
rect 278688 409566 278740 409572
rect 278700 408513 278728 409566
rect 278686 408504 278742 408513
rect 278686 408439 278742 408448
rect 281078 406600 281134 406609
rect 281078 406535 281134 406544
rect 278596 406292 278648 406298
rect 278596 406234 278648 406240
rect 277308 406224 277360 406230
rect 277308 406166 277360 406172
rect 275928 406156 275980 406162
rect 275928 406098 275980 406104
rect 243728 405884 243780 405890
rect 243728 405826 243780 405832
rect 281092 405822 281120 406535
rect 281460 406366 281488 572698
rect 282840 407114 282868 572698
rect 284220 412634 284248 572698
rect 284128 412606 284248 412634
rect 282828 407108 282880 407114
rect 282828 407050 282880 407056
rect 284128 407046 284156 412606
rect 284208 408332 284260 408338
rect 284208 408274 284260 408280
rect 284220 407153 284248 408274
rect 284206 407144 284262 407153
rect 284206 407079 284262 407088
rect 284116 407040 284168 407046
rect 284116 406982 284168 406988
rect 285600 406978 285628 575878
rect 286508 408604 286560 408610
rect 286508 408546 286560 408552
rect 286520 408377 286548 408546
rect 286506 408368 286562 408377
rect 286506 408303 286562 408312
rect 285588 406972 285640 406978
rect 285588 406914 285640 406920
rect 286980 406910 287008 575878
rect 288314 575634 288342 575892
rect 288314 575606 288388 575634
rect 286968 406904 287020 406910
rect 286968 406846 287020 406852
rect 288360 406842 288388 575606
rect 300768 407244 300820 407250
rect 300768 407186 300820 407192
rect 299388 407176 299440 407182
rect 299386 407144 299388 407153
rect 300780 407153 300808 407186
rect 299440 407144 299442 407153
rect 299386 407079 299442 407088
rect 300766 407144 300822 407153
rect 300766 407079 300822 407088
rect 288348 406836 288400 406842
rect 288348 406778 288400 406784
rect 281448 406360 281500 406366
rect 281448 406302 281500 406308
rect 281080 405816 281132 405822
rect 281080 405758 281132 405764
rect 316696 400994 316724 679254
rect 316776 679040 316828 679046
rect 316776 678982 316828 678988
rect 316684 400988 316736 400994
rect 316684 400930 316736 400936
rect 316788 400926 316816 678982
rect 323676 670744 323728 670750
rect 323676 670686 323728 670692
rect 320824 627972 320876 627978
rect 320824 627914 320876 627920
rect 320836 623082 320864 627914
rect 320824 623076 320876 623082
rect 320824 623018 320876 623024
rect 322204 572960 322256 572966
rect 322204 572902 322256 572908
rect 320916 501016 320968 501022
rect 320916 500958 320968 500964
rect 319536 409692 319588 409698
rect 319536 409634 319588 409640
rect 319444 408604 319496 408610
rect 319444 408546 319496 408552
rect 318248 408400 318300 408406
rect 318248 408342 318300 408348
rect 318062 407824 318118 407833
rect 318062 407759 318118 407768
rect 317604 407244 317656 407250
rect 317604 407186 317656 407192
rect 317512 407176 317564 407182
rect 317418 407144 317474 407153
rect 317512 407118 317564 407124
rect 317418 407079 317474 407088
rect 316866 406056 316922 406065
rect 316866 405991 316922 406000
rect 316776 400920 316828 400926
rect 316776 400862 316828 400868
rect 316880 389162 316908 405991
rect 316868 389156 316920 389162
rect 316868 389098 316920 389104
rect 278688 322244 278740 322250
rect 278688 322186 278740 322192
rect 223486 322008 223542 322017
rect 223486 321943 223542 321952
rect 228638 322008 228694 322017
rect 228638 321943 228694 321952
rect 179786 321872 179842 321881
rect 179512 321836 179564 321842
rect 223500 321842 223528 321943
rect 179786 321807 179842 321816
rect 223488 321836 223540 321842
rect 179512 321778 179564 321784
rect 179420 321768 179472 321774
rect 179418 321736 179420 321745
rect 179472 321736 179474 321745
rect 179418 321671 179474 321680
rect 179524 321609 179552 321778
rect 179800 321706 179828 321807
rect 223488 321778 223540 321784
rect 226340 321768 226392 321774
rect 226338 321736 226340 321745
rect 226392 321736 226394 321745
rect 179788 321700 179840 321706
rect 228652 321706 228680 321943
rect 226338 321671 226394 321680
rect 228640 321700 228692 321706
rect 179788 321642 179840 321648
rect 228640 321642 228692 321648
rect 229008 321700 229060 321706
rect 229008 321642 229060 321648
rect 204352 321632 204404 321638
rect 179510 321600 179566 321609
rect 204352 321574 204404 321580
rect 179510 321535 179566 321544
rect 180064 321564 180116 321570
rect 180064 321506 180116 321512
rect 178958 321464 179014 321473
rect 178958 321399 179014 321408
rect 179328 321428 179380 321434
rect 178592 321292 178644 321298
rect 178592 321234 178644 321240
rect 178604 320249 178632 321234
rect 178776 320476 178828 320482
rect 178776 320418 178828 320424
rect 178788 320249 178816 320418
rect 178590 320240 178646 320249
rect 178590 320175 178646 320184
rect 178774 320240 178830 320249
rect 178774 320175 178830 320184
rect 178500 319728 178552 319734
rect 178500 319670 178552 319676
rect 178408 311840 178460 311846
rect 178408 311782 178460 311788
rect 178316 296880 178368 296886
rect 178316 296822 178368 296828
rect 178132 294024 178184 294030
rect 178132 293966 178184 293972
rect 178144 292574 178172 293966
rect 178144 292546 178264 292574
rect 178132 289876 178184 289882
rect 178132 289818 178184 289824
rect 178040 288992 178092 288998
rect 178040 288934 178092 288940
rect 178052 205766 178080 288934
rect 178040 205760 178092 205766
rect 178040 205702 178092 205708
rect 178040 205624 178092 205630
rect 178040 205566 178092 205572
rect 177948 202972 178000 202978
rect 177948 202914 178000 202920
rect 176568 200524 176620 200530
rect 176568 200466 176620 200472
rect 178052 200326 178080 205566
rect 178144 200666 178172 289818
rect 178132 200660 178184 200666
rect 178132 200602 178184 200608
rect 178236 200598 178264 292546
rect 178328 210594 178356 296822
rect 178408 296812 178460 296818
rect 178408 296754 178460 296760
rect 178316 210588 178368 210594
rect 178316 210530 178368 210536
rect 178420 210474 178448 296754
rect 178328 210446 178448 210474
rect 178224 200592 178276 200598
rect 178224 200534 178276 200540
rect 178328 200394 178356 210446
rect 178408 210384 178460 210390
rect 178408 210326 178460 210332
rect 178420 205970 178448 210326
rect 178512 205970 178540 319670
rect 178592 319524 178644 319530
rect 178592 319466 178644 319472
rect 178604 205970 178632 319466
rect 178868 319388 178920 319394
rect 178868 319330 178920 319336
rect 178776 319320 178828 319326
rect 178776 319262 178828 319268
rect 178684 319184 178736 319190
rect 178684 319126 178736 319132
rect 178696 283082 178724 319126
rect 178684 283076 178736 283082
rect 178684 283018 178736 283024
rect 178684 282940 178736 282946
rect 178684 282882 178736 282888
rect 178696 267753 178724 282882
rect 178682 267744 178738 267753
rect 178682 267679 178738 267688
rect 178684 267640 178736 267646
rect 178684 267582 178736 267588
rect 178696 258126 178724 267582
rect 178684 258120 178736 258126
rect 178684 258062 178736 258068
rect 178684 257984 178736 257990
rect 178684 257926 178736 257932
rect 178408 205964 178460 205970
rect 178408 205906 178460 205912
rect 178500 205964 178552 205970
rect 178500 205906 178552 205912
rect 178592 205964 178644 205970
rect 178592 205906 178644 205912
rect 178696 205873 178724 257926
rect 178406 205864 178462 205873
rect 178406 205799 178462 205808
rect 178682 205864 178738 205873
rect 178682 205799 178738 205808
rect 178420 200462 178448 205799
rect 178500 205692 178552 205698
rect 178500 205634 178552 205640
rect 178592 205692 178644 205698
rect 178592 205634 178644 205640
rect 178684 205692 178736 205698
rect 178684 205634 178736 205640
rect 178512 203250 178540 205634
rect 178500 203244 178552 203250
rect 178500 203186 178552 203192
rect 178500 203108 178552 203114
rect 178500 203050 178552 203056
rect 178408 200456 178460 200462
rect 178408 200398 178460 200404
rect 178316 200388 178368 200394
rect 178316 200330 178368 200336
rect 178040 200320 178092 200326
rect 178040 200262 178092 200268
rect 178512 200258 178540 203050
rect 178604 201006 178632 205634
rect 178592 201000 178644 201006
rect 178592 200942 178644 200948
rect 178500 200252 178552 200258
rect 178500 200194 178552 200200
rect 178696 200190 178724 205634
rect 178788 200734 178816 319262
rect 178880 200870 178908 319330
rect 178868 200864 178920 200870
rect 178868 200806 178920 200812
rect 178776 200728 178828 200734
rect 178776 200670 178828 200676
rect 178972 200433 179000 321399
rect 179328 321370 179380 321376
rect 179144 321360 179196 321366
rect 179144 321302 179196 321308
rect 179052 320544 179104 320550
rect 179052 320486 179104 320492
rect 179064 201074 179092 320486
rect 179156 201210 179184 321302
rect 179236 320816 179288 320822
rect 179236 320758 179288 320764
rect 179248 210594 179276 320758
rect 179236 210588 179288 210594
rect 179236 210530 179288 210536
rect 179340 210474 179368 321370
rect 179510 321192 179566 321201
rect 179510 321127 179566 321136
rect 179524 320618 179552 321127
rect 179420 320612 179472 320618
rect 179420 320554 179472 320560
rect 179512 320612 179564 320618
rect 179512 320554 179564 320560
rect 179432 320346 179460 320554
rect 179420 320340 179472 320346
rect 179420 320282 179472 320288
rect 179524 320249 179552 320554
rect 179972 320408 180024 320414
rect 179972 320350 180024 320356
rect 179880 320340 179932 320346
rect 179880 320282 179932 320288
rect 179510 320240 179566 320249
rect 179510 320175 179566 320184
rect 179788 320068 179840 320074
rect 179788 320010 179840 320016
rect 179696 319932 179748 319938
rect 179696 319874 179748 319880
rect 179604 319796 179656 319802
rect 179604 319738 179656 319744
rect 179420 319660 179472 319666
rect 179420 319602 179472 319608
rect 179432 319462 179460 319602
rect 179512 319592 179564 319598
rect 179512 319534 179564 319540
rect 179420 319456 179472 319462
rect 179420 319398 179472 319404
rect 179420 319252 179472 319258
rect 179420 319194 179472 319200
rect 179432 215354 179460 319194
rect 179420 215348 179472 215354
rect 179420 215290 179472 215296
rect 179420 215212 179472 215218
rect 179420 215154 179472 215160
rect 179432 210730 179460 215154
rect 179420 210724 179472 210730
rect 179420 210666 179472 210672
rect 179420 210588 179472 210594
rect 179420 210530 179472 210536
rect 179248 210446 179368 210474
rect 179144 201204 179196 201210
rect 179144 201146 179196 201152
rect 179248 201142 179276 210446
rect 179328 210384 179380 210390
rect 179328 210326 179380 210332
rect 179340 205970 179368 210326
rect 179328 205964 179380 205970
rect 179328 205906 179380 205912
rect 179326 205864 179382 205873
rect 179326 205799 179382 205808
rect 179340 203833 179368 205799
rect 179326 203824 179382 203833
rect 179326 203759 179382 203768
rect 179432 203114 179460 210530
rect 179524 203454 179552 319534
rect 179616 319462 179644 319738
rect 179604 319456 179656 319462
rect 179604 319398 179656 319404
rect 179616 318458 179644 319398
rect 179708 319394 179736 319874
rect 179696 319388 179748 319394
rect 179696 319330 179748 319336
rect 179708 318594 179736 319330
rect 179800 319258 179828 320010
rect 179788 319252 179840 319258
rect 179788 319194 179840 319200
rect 179708 318566 179828 318594
rect 179616 318430 179736 318458
rect 179604 318368 179656 318374
rect 179604 318310 179656 318316
rect 179616 258092 179644 318310
rect 179604 258086 179656 258092
rect 179604 258028 179656 258034
rect 179708 257938 179736 318430
rect 179800 318374 179828 318566
rect 179788 318368 179840 318374
rect 179788 318310 179840 318316
rect 179892 318186 179920 320282
rect 179616 257910 179736 257938
rect 179800 318158 179920 318186
rect 179616 244050 179644 257910
rect 179696 257848 179748 257854
rect 179696 257790 179748 257796
rect 179708 253910 179736 257790
rect 179696 253904 179748 253910
rect 179696 253846 179748 253852
rect 179696 253768 179748 253774
rect 179696 253710 179748 253716
rect 179708 244390 179736 253710
rect 179696 244384 179748 244390
rect 179696 244326 179748 244332
rect 179696 244180 179748 244186
rect 179696 244122 179748 244128
rect 179604 244044 179656 244050
rect 179604 243986 179656 243992
rect 179602 243944 179658 243953
rect 179602 243879 179658 243888
rect 179616 236473 179644 243879
rect 179602 236464 179658 236473
rect 179602 236399 179658 236408
rect 179708 234734 179736 244122
rect 179604 234728 179656 234734
rect 179604 234670 179656 234676
rect 179696 234728 179748 234734
rect 179696 234670 179748 234676
rect 179616 225078 179644 234670
rect 179696 234626 179748 234632
rect 179696 234568 179748 234574
rect 179604 225072 179656 225078
rect 179604 225014 179656 225020
rect 179604 224868 179656 224874
rect 179604 224810 179656 224816
rect 179616 210594 179644 224810
rect 179604 210588 179656 210594
rect 179604 210530 179656 210536
rect 179708 210474 179736 234568
rect 179616 210446 179736 210474
rect 179512 203448 179564 203454
rect 179512 203390 179564 203396
rect 179616 203182 179644 210446
rect 179696 210384 179748 210390
rect 179696 210326 179748 210332
rect 179708 205834 179736 210326
rect 179696 205828 179748 205834
rect 179696 205770 179748 205776
rect 179696 205692 179748 205698
rect 179696 205634 179748 205640
rect 179604 203176 179656 203182
rect 179604 203118 179656 203124
rect 179420 203108 179472 203114
rect 179420 203050 179472 203056
rect 179708 203046 179736 205634
rect 179696 203040 179748 203046
rect 179696 202982 179748 202988
rect 179800 201482 179828 318158
rect 179984 318050 180012 320350
rect 179892 318022 180012 318050
rect 179788 201476 179840 201482
rect 179788 201418 179840 201424
rect 179892 201414 179920 318022
rect 180076 316034 180104 321506
rect 180154 321464 180210 321473
rect 180154 321399 180210 321408
rect 180168 320210 180196 321399
rect 203156 321292 203208 321298
rect 203156 321234 203208 321240
rect 202788 320340 202840 320346
rect 202788 320282 202840 320288
rect 180156 320204 180208 320210
rect 180156 320146 180208 320152
rect 200764 320136 200816 320142
rect 200762 320104 200764 320113
rect 200816 320104 200818 320113
rect 200762 320039 200818 320048
rect 180524 319660 180576 319666
rect 180524 319602 180576 319608
rect 180536 318889 180564 319602
rect 196070 319424 196126 319433
rect 196070 319359 196126 319368
rect 197358 319424 197414 319433
rect 197358 319359 197414 319368
rect 198738 319424 198794 319433
rect 198738 319359 198794 319368
rect 196084 319122 196112 319359
rect 196072 319116 196124 319122
rect 196072 319058 196124 319064
rect 195992 318918 196020 318949
rect 195980 318912 196032 318918
rect 180522 318880 180578 318889
rect 180522 318815 180578 318824
rect 195978 318880 195980 318889
rect 196032 318880 196034 318889
rect 195978 318815 196034 318824
rect 179984 316006 180104 316034
rect 179880 201408 179932 201414
rect 179880 201350 179932 201356
rect 179984 201346 180012 316006
rect 195992 291242 196020 318815
rect 195980 291236 196032 291242
rect 195980 291178 196032 291184
rect 196084 291122 196112 319058
rect 197372 319054 197400 319359
rect 197360 319048 197412 319054
rect 197360 318990 197412 318996
rect 197372 296886 197400 318990
rect 198752 318986 198780 319359
rect 198740 318980 198792 318986
rect 198740 318922 198792 318928
rect 197360 296880 197412 296886
rect 197360 296822 197412 296828
rect 197372 296682 197400 296822
rect 198752 296818 198780 318922
rect 200776 298110 200804 320039
rect 201498 319288 201554 319297
rect 201498 319223 201554 319232
rect 201512 319190 201540 319223
rect 202800 319190 202828 320282
rect 203168 320113 203196 321234
rect 204364 320113 204392 321574
rect 219438 321464 219494 321473
rect 219438 321399 219440 321408
rect 219492 321399 219494 321408
rect 220450 321464 220506 321473
rect 220450 321399 220506 321408
rect 220636 321428 220688 321434
rect 219440 321370 219492 321376
rect 220464 321366 220492 321399
rect 220636 321370 220688 321376
rect 220452 321360 220504 321366
rect 220452 321302 220504 321308
rect 211068 320816 211120 320822
rect 211068 320758 211120 320764
rect 207294 320648 207350 320657
rect 207294 320583 207350 320592
rect 204904 320272 204956 320278
rect 204904 320214 204956 320220
rect 204916 320142 204944 320214
rect 204904 320136 204956 320142
rect 203154 320104 203210 320113
rect 203154 320039 203210 320048
rect 203798 320104 203854 320113
rect 203798 320039 203854 320048
rect 204350 320104 204406 320113
rect 204904 320078 204956 320084
rect 204350 320039 204406 320048
rect 201500 319184 201552 319190
rect 201500 319126 201552 319132
rect 202144 319184 202196 319190
rect 202144 319126 202196 319132
rect 202788 319184 202840 319190
rect 202788 319126 202840 319132
rect 200764 298104 200816 298110
rect 200764 298046 200816 298052
rect 202156 298042 202184 319126
rect 203812 318374 203840 320039
rect 204258 319152 204314 319161
rect 204258 319087 204314 319096
rect 204272 318850 204300 319087
rect 204260 318844 204312 318850
rect 204260 318786 204312 318792
rect 203800 318368 203852 318374
rect 203800 318310 203852 318316
rect 202144 298036 202196 298042
rect 202144 297978 202196 297984
rect 198740 296812 198792 296818
rect 198740 296754 198792 296760
rect 197360 296676 197412 296682
rect 197360 296618 197412 296624
rect 198752 296614 198780 296754
rect 198740 296608 198792 296614
rect 198740 296550 198792 296556
rect 196164 291236 196216 291242
rect 196164 291178 196216 291184
rect 195992 291094 196112 291122
rect 195992 289066 196020 291094
rect 196176 290986 196204 291178
rect 196084 290958 196204 290986
rect 180708 289060 180760 289066
rect 180708 289002 180760 289008
rect 195980 289060 196032 289066
rect 195980 289002 196032 289008
rect 180338 287464 180394 287473
rect 180720 287434 180748 289002
rect 195992 287774 196020 289002
rect 196084 288998 196112 290958
rect 204272 289882 204300 318786
rect 204364 294030 204392 320039
rect 207308 319734 207336 320583
rect 208400 320204 208452 320210
rect 208400 320146 208452 320152
rect 208412 319734 208440 320146
rect 211080 319870 211108 320758
rect 215116 320612 215168 320618
rect 215116 320554 215168 320560
rect 211802 320104 211858 320113
rect 211802 320039 211858 320048
rect 211816 320006 211844 320039
rect 211804 320000 211856 320006
rect 215128 319977 215156 320554
rect 216404 320544 216456 320550
rect 216404 320486 216456 320492
rect 211804 319942 211856 319948
rect 215114 319968 215170 319977
rect 211068 319864 211120 319870
rect 210422 319832 210478 319841
rect 211068 319806 211120 319812
rect 210422 319767 210424 319776
rect 210476 319767 210478 319776
rect 210424 319738 210476 319744
rect 207296 319728 207348 319734
rect 207296 319670 207348 319676
rect 208400 319728 208452 319734
rect 208400 319670 208452 319676
rect 206282 319288 206338 319297
rect 206282 319223 206338 319232
rect 204352 294024 204404 294030
rect 204352 293966 204404 293972
rect 204364 293418 204392 293966
rect 204352 293412 204404 293418
rect 204352 293354 204404 293360
rect 206296 291854 206324 319223
rect 207308 318442 207336 319670
rect 209042 319288 209098 319297
rect 209042 319223 209098 319232
rect 207296 318436 207348 318442
rect 207296 318378 207348 318384
rect 206284 291848 206336 291854
rect 206284 291790 206336 291796
rect 204260 289876 204312 289882
rect 204260 289818 204312 289824
rect 204720 289876 204772 289882
rect 204720 289818 204772 289824
rect 204732 289338 204760 289818
rect 204720 289332 204772 289338
rect 204720 289274 204772 289280
rect 196072 288992 196124 288998
rect 196072 288934 196124 288940
rect 195980 287768 196032 287774
rect 195980 287710 196032 287716
rect 196084 287706 196112 288934
rect 209056 287910 209084 319223
rect 209320 298172 209372 298178
rect 209320 298114 209372 298120
rect 209332 291145 209360 298114
rect 209318 291136 209374 291145
rect 209318 291071 209374 291080
rect 209044 287904 209096 287910
rect 209044 287846 209096 287852
rect 210436 287842 210464 319738
rect 211342 319152 211398 319161
rect 211342 319087 211344 319096
rect 211396 319087 211398 319096
rect 211344 319058 211396 319064
rect 211068 300892 211120 300898
rect 211068 300834 211120 300840
rect 211080 291145 211108 300834
rect 211066 291136 211122 291145
rect 211066 291071 211122 291080
rect 211816 287978 211844 319942
rect 215114 319903 215170 319912
rect 213184 319592 213236 319598
rect 213184 319534 213236 319540
rect 213196 319433 213224 319534
rect 213182 319424 213238 319433
rect 213182 319359 213238 319368
rect 211986 319152 212042 319161
rect 211986 319087 212042 319096
rect 212000 288046 212028 319087
rect 213196 293350 213224 319359
rect 213828 303680 213880 303686
rect 213828 303622 213880 303628
rect 213184 293344 213236 293350
rect 213184 293286 213236 293292
rect 213840 291145 213868 303622
rect 213826 291136 213882 291145
rect 213826 291071 213882 291080
rect 215128 289474 215156 319903
rect 216416 319705 216444 320486
rect 216680 320476 216732 320482
rect 216680 320418 216732 320424
rect 216692 319705 216720 320418
rect 218060 320408 218112 320414
rect 218060 320350 218112 320356
rect 218072 319705 218100 320350
rect 216402 319696 216458 319705
rect 216402 319631 216458 319640
rect 216678 319696 216734 319705
rect 216678 319631 216734 319640
rect 217874 319696 217930 319705
rect 217874 319631 217930 319640
rect 218058 319696 218114 319705
rect 218058 319631 218114 319640
rect 219254 319696 219310 319705
rect 219254 319631 219310 319640
rect 216416 292126 216444 319631
rect 216496 306400 216548 306406
rect 216496 306342 216548 306348
rect 216404 292120 216456 292126
rect 216404 292062 216456 292068
rect 216508 291145 216536 306342
rect 216494 291136 216550 291145
rect 216494 291071 216550 291080
rect 215116 289468 215168 289474
rect 215116 289410 215168 289416
rect 217888 289406 217916 319631
rect 219268 312594 219296 319631
rect 219256 312588 219308 312594
rect 219256 312530 219308 312536
rect 219348 309188 219400 309194
rect 219348 309130 219400 309136
rect 219360 291145 219388 309130
rect 220464 292194 220492 321302
rect 220648 294642 220676 321370
rect 221830 320648 221886 320657
rect 221830 320583 221886 320592
rect 221844 319870 221872 320583
rect 224144 320142 224172 320173
rect 224132 320136 224184 320142
rect 224130 320104 224132 320113
rect 224184 320104 224186 320113
rect 224130 320039 224186 320048
rect 227534 320104 227590 320113
rect 227534 320039 227590 320048
rect 221832 319864 221884 319870
rect 221832 319806 221884 319812
rect 222108 319864 222160 319870
rect 222108 319806 222160 319812
rect 222120 318510 222148 319806
rect 222844 319728 222896 319734
rect 222844 319670 222896 319676
rect 222856 319433 222884 319670
rect 222842 319424 222898 319433
rect 222842 319359 222898 319368
rect 222108 318504 222160 318510
rect 222108 318446 222160 318452
rect 222108 311908 222160 311914
rect 222108 311850 222160 311856
rect 220636 294636 220688 294642
rect 220636 294578 220688 294584
rect 220452 292188 220504 292194
rect 220452 292130 220504 292136
rect 222120 291145 222148 311850
rect 219346 291136 219402 291145
rect 219346 291071 219402 291080
rect 222106 291136 222162 291145
rect 222106 291071 222162 291080
rect 222856 289542 222884 319359
rect 224144 318918 224172 320039
rect 226982 319968 227038 319977
rect 226982 319903 227038 319912
rect 225602 319288 225658 319297
rect 225602 319223 225658 319232
rect 225616 319190 225644 319223
rect 225604 319184 225656 319190
rect 225604 319126 225656 319132
rect 224132 318912 224184 318918
rect 224132 318854 224184 318860
rect 223488 314764 223540 314770
rect 223488 314706 223540 314712
rect 223500 291145 223528 314706
rect 223486 291136 223542 291145
rect 223486 291071 223542 291080
rect 222844 289536 222896 289542
rect 222844 289478 222896 289484
rect 217876 289400 217928 289406
rect 217876 289342 217928 289348
rect 225616 288386 225644 319126
rect 226248 316056 226300 316062
rect 226248 315998 226300 316004
rect 226260 291145 226288 315998
rect 226246 291136 226302 291145
rect 226246 291071 226302 291080
rect 225604 288380 225656 288386
rect 225604 288322 225656 288328
rect 226996 288318 227024 319903
rect 226984 288312 227036 288318
rect 226984 288254 227036 288260
rect 227548 288250 227576 320039
rect 228916 318844 228968 318850
rect 228916 318786 228968 318792
rect 228928 291145 228956 318786
rect 228914 291136 228970 291145
rect 228914 291071 228970 291080
rect 229020 289814 229048 321642
rect 231768 321632 231820 321638
rect 231768 321574 231820 321580
rect 231214 320104 231270 320113
rect 231214 320039 231270 320048
rect 229558 319968 229614 319977
rect 229558 319903 229560 319912
rect 229612 319903 229614 319912
rect 229560 319874 229612 319880
rect 229572 316034 229600 319874
rect 231228 319530 231256 320039
rect 231216 319524 231268 319530
rect 231216 319466 231268 319472
rect 231676 319524 231728 319530
rect 231676 319466 231728 319472
rect 231688 318986 231716 319466
rect 231676 318980 231728 318986
rect 231676 318922 231728 318928
rect 229572 316006 229784 316034
rect 229008 289808 229060 289814
rect 229008 289750 229060 289756
rect 229756 289746 229784 316006
rect 231780 291145 231808 321574
rect 246948 321428 247000 321434
rect 246948 321370 247000 321376
rect 241428 321292 241480 321298
rect 241428 321234 241480 321240
rect 232044 320748 232096 320754
rect 232044 320690 232096 320696
rect 231858 319696 231914 319705
rect 231858 319631 231860 319640
rect 231912 319631 231914 319640
rect 231860 319602 231912 319608
rect 232056 319530 232084 320690
rect 233884 320680 233936 320686
rect 233884 320622 233936 320628
rect 232502 319696 232558 319705
rect 232502 319631 232558 319640
rect 232044 319524 232096 319530
rect 232044 319466 232096 319472
rect 231766 291136 231822 291145
rect 231766 291071 231822 291080
rect 232516 290358 232544 319631
rect 233896 319598 233924 320622
rect 236644 320068 236696 320074
rect 236644 320010 236696 320016
rect 233884 319592 233936 319598
rect 236656 319569 236684 320010
rect 233884 319534 233936 319540
rect 236642 319560 236698 319569
rect 236642 319495 236698 319504
rect 233884 319456 233936 319462
rect 233884 319398 233936 319404
rect 233896 318889 233924 319398
rect 234068 319388 234120 319394
rect 234068 319330 234120 319336
rect 234080 319297 234108 319330
rect 235276 319326 235304 319357
rect 235264 319320 235316 319326
rect 234066 319288 234122 319297
rect 234066 319223 234122 319232
rect 235262 319288 235264 319297
rect 235316 319288 235318 319297
rect 235262 319223 235318 319232
rect 233882 318880 233938 318889
rect 233882 318815 233938 318824
rect 233896 292466 233924 318815
rect 234080 292534 234108 319223
rect 235276 293894 235304 319223
rect 235264 293888 235316 293894
rect 235264 293830 235316 293836
rect 236656 293826 236684 319495
rect 238024 319252 238076 319258
rect 238024 319194 238076 319200
rect 238036 319161 238064 319194
rect 238022 319152 238078 319161
rect 238022 319087 238078 319096
rect 238036 295322 238064 319087
rect 239402 319016 239458 319025
rect 239402 318951 239458 318960
rect 238668 315308 238720 315314
rect 238668 315250 238720 315256
rect 238024 295316 238076 295322
rect 238024 295258 238076 295264
rect 236644 293820 236696 293826
rect 236644 293762 236696 293768
rect 234068 292528 234120 292534
rect 234068 292470 234120 292476
rect 233884 292460 233936 292466
rect 233884 292402 233936 292408
rect 237288 292256 237340 292262
rect 237288 292198 237340 292204
rect 237300 291009 237328 292198
rect 238680 291145 238708 315250
rect 239416 294710 239444 318951
rect 239404 294704 239456 294710
rect 239404 294646 239456 294652
rect 241440 291145 241468 321234
rect 244188 292324 244240 292330
rect 244188 292266 244240 292272
rect 244200 291145 244228 292266
rect 246960 291145 246988 321370
rect 253848 321360 253900 321366
rect 253848 321302 253900 321308
rect 251088 318640 251140 318646
rect 251088 318582 251140 318588
rect 249708 318572 249760 318578
rect 249708 318514 249760 318520
rect 249720 291145 249748 318514
rect 251100 291145 251128 318582
rect 253860 291145 253888 321302
rect 271788 319932 271840 319938
rect 271788 319874 271840 319880
rect 269028 319796 269080 319802
rect 269028 319738 269080 319744
rect 264888 319660 264940 319666
rect 264888 319602 264940 319608
rect 256608 319456 256660 319462
rect 256608 319398 256660 319404
rect 256620 291145 256648 319398
rect 259368 318708 259420 318714
rect 259368 318650 259420 318656
rect 259380 291145 259408 318650
rect 262128 292392 262180 292398
rect 262128 292334 262180 292340
rect 238666 291136 238722 291145
rect 238666 291071 238722 291080
rect 241426 291136 241482 291145
rect 241426 291071 241482 291080
rect 244186 291136 244242 291145
rect 244186 291071 244242 291080
rect 246946 291136 247002 291145
rect 246946 291071 247002 291080
rect 249706 291136 249762 291145
rect 249706 291071 249762 291080
rect 251086 291136 251142 291145
rect 251086 291071 251142 291080
rect 253846 291136 253902 291145
rect 253846 291071 253902 291080
rect 256606 291136 256662 291145
rect 256606 291071 256662 291080
rect 259366 291136 259422 291145
rect 259366 291071 259422 291080
rect 237286 291000 237342 291009
rect 237286 290935 237342 290944
rect 262140 290465 262168 292334
rect 264900 291145 264928 319602
rect 266268 293480 266320 293486
rect 266268 293422 266320 293428
rect 264886 291136 264942 291145
rect 264886 291071 264942 291080
rect 266280 290737 266308 293422
rect 269040 291145 269068 319738
rect 271800 291145 271828 319874
rect 277308 319864 277360 319870
rect 277308 319806 277360 319812
rect 274548 319728 274600 319734
rect 274548 319670 274600 319676
rect 274560 291145 274588 319670
rect 277320 291145 277348 319806
rect 269026 291136 269082 291145
rect 269026 291071 269082 291080
rect 271786 291136 271842 291145
rect 271786 291071 271842 291080
rect 274546 291136 274602 291145
rect 274546 291071 274602 291080
rect 277306 291136 277362 291145
rect 277306 291071 277362 291080
rect 278700 290737 278728 322186
rect 303068 319592 303120 319598
rect 303068 319534 303120 319540
rect 302884 319524 302936 319530
rect 302884 319466 302936 319472
rect 302896 319297 302924 319466
rect 303080 319433 303108 319534
rect 303066 319424 303122 319433
rect 303066 319359 303122 319368
rect 302882 319288 302938 319297
rect 302882 319223 302938 319232
rect 281448 318776 281500 318782
rect 281448 318718 281500 318724
rect 281460 291145 281488 318718
rect 284208 291780 284260 291786
rect 284208 291722 284260 291728
rect 284220 291145 284248 291722
rect 281446 291136 281502 291145
rect 281446 291071 281502 291080
rect 284206 291136 284262 291145
rect 284206 291071 284262 291080
rect 266266 290728 266322 290737
rect 266266 290663 266322 290672
rect 278686 290728 278742 290737
rect 278686 290663 278742 290672
rect 299664 290556 299716 290562
rect 299664 290498 299716 290504
rect 262126 290456 262182 290465
rect 262126 290391 262182 290400
rect 299020 290420 299072 290426
rect 299020 290362 299072 290368
rect 232504 290352 232556 290358
rect 232504 290294 232556 290300
rect 234528 290284 234580 290290
rect 234528 290226 234580 290232
rect 234540 290057 234568 290226
rect 286600 290216 286652 290222
rect 286600 290158 286652 290164
rect 234526 290048 234582 290057
rect 234526 289983 234582 289992
rect 286612 289921 286640 290158
rect 299032 289921 299060 290362
rect 299676 289921 299704 290498
rect 286598 289912 286654 289921
rect 286598 289847 286654 289856
rect 299018 289912 299074 289921
rect 299018 289847 299074 289856
rect 299662 289912 299718 289921
rect 299662 289847 299718 289856
rect 229744 289740 229796 289746
rect 229744 289682 229796 289688
rect 299032 289678 299060 289847
rect 299020 289672 299072 289678
rect 299020 289614 299072 289620
rect 302896 289610 302924 319223
rect 303080 293554 303108 319359
rect 316776 318980 316828 318986
rect 316776 318922 316828 318928
rect 316684 318912 316736 318918
rect 316684 318854 316736 318860
rect 316500 294704 316552 294710
rect 316500 294646 316552 294652
rect 316512 294030 316540 294646
rect 316500 294024 316552 294030
rect 316500 293966 316552 293972
rect 303068 293548 303120 293554
rect 303068 293490 303120 293496
rect 316512 291938 316540 293966
rect 316512 291910 316632 291938
rect 310796 290420 310848 290426
rect 310796 290362 310848 290368
rect 310808 289921 310836 290362
rect 310794 289912 310850 289921
rect 310794 289847 310850 289856
rect 302884 289604 302936 289610
rect 302884 289546 302936 289552
rect 227536 288244 227588 288250
rect 227536 288186 227588 288192
rect 211988 288040 212040 288046
rect 211988 287982 212040 287988
rect 211804 287972 211856 287978
rect 211804 287914 211856 287920
rect 210424 287836 210476 287842
rect 210424 287778 210476 287784
rect 196072 287700 196124 287706
rect 196072 287642 196124 287648
rect 180338 287399 180340 287408
rect 180392 287399 180394 287408
rect 180708 287428 180760 287434
rect 180340 287370 180392 287376
rect 180708 287370 180760 287376
rect 229742 203552 229798 203561
rect 229742 203487 229798 203496
rect 231122 203552 231178 203561
rect 231122 203487 231178 203496
rect 232226 203552 232282 203561
rect 232226 203487 232282 203496
rect 233330 203552 233386 203561
rect 233330 203487 233386 203496
rect 234434 203552 234490 203561
rect 234434 203487 234490 203496
rect 235722 203552 235778 203561
rect 235722 203487 235778 203496
rect 237010 203552 237066 203561
rect 237010 203487 237066 203496
rect 238022 203552 238078 203561
rect 238022 203487 238078 203496
rect 229756 203318 229784 203487
rect 231136 203386 231164 203487
rect 231124 203380 231176 203386
rect 231124 203322 231176 203328
rect 180064 203312 180116 203318
rect 180064 203254 180116 203260
rect 229744 203312 229796 203318
rect 229744 203254 229796 203260
rect 179972 201340 180024 201346
rect 179972 201282 180024 201288
rect 180076 201278 180104 203254
rect 232240 203250 232268 203487
rect 232228 203244 232280 203250
rect 232228 203186 232280 203192
rect 233344 203182 233372 203487
rect 233332 203176 233384 203182
rect 233332 203118 233384 203124
rect 234448 203114 234476 203487
rect 234436 203108 234488 203114
rect 234436 203050 234488 203056
rect 235736 203046 235764 203487
rect 235724 203040 235776 203046
rect 235724 202982 235776 202988
rect 237024 202910 237052 203487
rect 238036 202978 238064 203487
rect 238024 202972 238076 202978
rect 238024 202914 238076 202920
rect 237012 202904 237064 202910
rect 237012 202846 237064 202852
rect 316604 201482 316632 291910
rect 316696 287026 316724 318854
rect 316788 290970 316816 318922
rect 316776 290964 316828 290970
rect 316776 290906 316828 290912
rect 317432 290426 317460 407079
rect 317420 290420 317472 290426
rect 317420 290362 317472 290368
rect 317524 289678 317552 407118
rect 317616 290562 317644 407186
rect 318076 345030 318104 407759
rect 318154 405920 318210 405929
rect 318154 405855 318210 405864
rect 318168 389094 318196 405855
rect 318156 389088 318208 389094
rect 318156 389030 318208 389036
rect 318156 376780 318208 376786
rect 318156 376722 318208 376728
rect 318064 345024 318116 345030
rect 318064 344966 318116 344972
rect 318168 290630 318196 376722
rect 318260 376718 318288 408342
rect 318432 408264 318484 408270
rect 318432 408206 318484 408212
rect 318340 405816 318392 405822
rect 318340 405758 318392 405764
rect 318248 376712 318300 376718
rect 318248 376654 318300 376660
rect 318352 375358 318380 405758
rect 318340 375352 318392 375358
rect 318340 375294 318392 375300
rect 318248 374060 318300 374066
rect 318248 374002 318300 374008
rect 318260 290698 318288 374002
rect 318444 371890 318472 408206
rect 318524 407584 318576 407590
rect 318524 407526 318576 407532
rect 318432 371884 318484 371890
rect 318432 371826 318484 371832
rect 318340 371272 318392 371278
rect 318340 371214 318392 371220
rect 318352 290766 318380 371214
rect 318432 369912 318484 369918
rect 318432 369854 318484 369860
rect 318444 290834 318472 369854
rect 318536 368490 318564 407526
rect 319456 380730 319484 408546
rect 319444 380724 319496 380730
rect 319444 380666 319496 380672
rect 319444 378208 319496 378214
rect 319444 378150 319496 378156
rect 318524 368484 318576 368490
rect 318524 368426 318576 368432
rect 318524 324352 318576 324358
rect 318524 324294 318576 324300
rect 318432 290828 318484 290834
rect 318432 290770 318484 290776
rect 318340 290760 318392 290766
rect 318340 290702 318392 290708
rect 318248 290692 318300 290698
rect 318248 290634 318300 290640
rect 318156 290624 318208 290630
rect 318156 290566 318208 290572
rect 317604 290556 317656 290562
rect 317604 290498 317656 290504
rect 318536 290290 318564 324294
rect 318616 290556 318668 290562
rect 318616 290498 318668 290504
rect 318524 290284 318576 290290
rect 318524 290226 318576 290232
rect 317512 289672 317564 289678
rect 317512 289614 317564 289620
rect 318156 289604 318208 289610
rect 318156 289546 318208 289552
rect 317420 289536 317472 289542
rect 317420 289478 317472 289484
rect 316684 287020 316736 287026
rect 316684 286962 316736 286968
rect 317432 286958 317460 289478
rect 318064 287360 318116 287366
rect 318064 287302 318116 287308
rect 317420 286952 317472 286958
rect 317420 286894 317472 286900
rect 318076 273222 318104 287302
rect 318064 273216 318116 273222
rect 318064 273158 318116 273164
rect 318168 262886 318196 289546
rect 318156 262880 318208 262886
rect 318156 262822 318208 262828
rect 318628 259418 318656 290498
rect 318708 290420 318760 290426
rect 318708 290362 318760 290368
rect 318720 289134 318748 290362
rect 319456 290222 319484 378150
rect 319548 357406 319576 409634
rect 319628 408196 319680 408202
rect 319628 408138 319680 408144
rect 319640 359514 319668 408138
rect 320086 401704 320142 401713
rect 320086 401639 320088 401648
rect 320140 401639 320142 401648
rect 320088 401610 320140 401616
rect 320824 397520 320876 397526
rect 320824 397462 320876 397468
rect 319628 359508 319680 359514
rect 319628 359450 319680 359456
rect 319536 357400 319588 357406
rect 319536 357342 319588 357348
rect 319534 341728 319590 341737
rect 319534 341663 319590 341672
rect 319444 290216 319496 290222
rect 319444 290158 319496 290164
rect 318708 289128 318760 289134
rect 318708 289070 318760 289076
rect 319442 283248 319498 283257
rect 319442 283183 319498 283192
rect 319456 271862 319484 283183
rect 319444 271856 319496 271862
rect 319444 271798 319496 271804
rect 319444 262200 319496 262206
rect 319444 262142 319496 262148
rect 319456 261526 319484 262142
rect 319444 261520 319496 261526
rect 319444 261462 319496 261468
rect 318616 259412 318668 259418
rect 318616 259354 318668 259360
rect 318064 256216 318116 256222
rect 318064 256158 318116 256164
rect 317418 223408 317474 223417
rect 317418 223343 317474 223352
rect 317432 203930 317460 223343
rect 317510 221776 317566 221785
rect 317510 221711 317566 221720
rect 317420 203924 317472 203930
rect 317420 203866 317472 203872
rect 317524 203522 317552 221711
rect 317602 217696 317658 217705
rect 317602 217631 317658 217640
rect 317616 203998 317644 217631
rect 317604 203992 317656 203998
rect 317604 203934 317656 203940
rect 317512 203516 317564 203522
rect 317512 203458 317564 203464
rect 224960 201476 225012 201482
rect 224960 201418 225012 201424
rect 238944 201476 238996 201482
rect 238944 201418 238996 201424
rect 316592 201476 316644 201482
rect 316592 201418 316644 201424
rect 223580 201408 223632 201414
rect 195978 201376 196034 201385
rect 195978 201311 196034 201320
rect 196162 201376 196218 201385
rect 196162 201311 196218 201320
rect 197358 201376 197414 201385
rect 197358 201311 197414 201320
rect 198738 201376 198794 201385
rect 198738 201311 198794 201320
rect 200118 201376 200174 201385
rect 200118 201311 200174 201320
rect 204350 201376 204406 201385
rect 204350 201311 204406 201320
rect 211250 201376 211306 201385
rect 211250 201311 211306 201320
rect 219990 201376 220046 201385
rect 219990 201311 220046 201320
rect 222198 201376 222254 201385
rect 222198 201311 222200 201320
rect 195992 201278 196020 201311
rect 180064 201272 180116 201278
rect 180064 201214 180116 201220
rect 195980 201272 196032 201278
rect 195980 201214 196032 201220
rect 179236 201136 179288 201142
rect 179236 201078 179288 201084
rect 179052 201068 179104 201074
rect 179052 201010 179104 201016
rect 178958 200424 179014 200433
rect 178958 200359 179014 200368
rect 196176 200258 196204 201311
rect 197372 200326 197400 201311
rect 198752 200394 198780 201311
rect 200132 200530 200160 201311
rect 204258 201240 204314 201249
rect 204258 201175 204314 201184
rect 204272 200598 204300 201175
rect 204364 200666 204392 201311
rect 211158 201104 211214 201113
rect 211158 201039 211214 201048
rect 211172 201006 211200 201039
rect 211160 201000 211212 201006
rect 211160 200942 211212 200948
rect 211264 200870 211292 201311
rect 215298 201240 215354 201249
rect 215298 201175 215354 201184
rect 219438 201240 219494 201249
rect 220004 201210 220032 201311
rect 222252 201311 222254 201320
rect 223578 201376 223580 201385
rect 224972 201385 225000 201418
rect 238956 201385 238984 201418
rect 302240 201408 302292 201414
rect 223632 201376 223634 201385
rect 223578 201311 223634 201320
rect 224958 201376 225014 201385
rect 224958 201311 225014 201320
rect 238942 201376 238998 201385
rect 303160 201408 303212 201414
rect 302240 201350 302292 201356
rect 303158 201376 303160 201385
rect 303212 201376 303214 201385
rect 238942 201311 238998 201320
rect 222200 201282 222252 201288
rect 219438 201175 219494 201184
rect 219992 201204 220044 201210
rect 215312 201074 215340 201175
rect 219452 201142 219480 201175
rect 219992 201146 220044 201152
rect 219440 201136 219492 201142
rect 219440 201078 219492 201084
rect 215300 201068 215352 201074
rect 215300 201010 215352 201016
rect 302252 200938 302280 201350
rect 302332 201340 302384 201346
rect 303158 201311 303214 201320
rect 303526 201376 303582 201385
rect 303526 201311 303528 201320
rect 302332 201282 302384 201288
rect 303580 201311 303582 201320
rect 303528 201282 303580 201288
rect 302240 200932 302292 200938
rect 302240 200874 302292 200880
rect 211252 200864 211304 200870
rect 209870 200832 209926 200841
rect 211252 200806 211304 200812
rect 302344 200802 302372 201282
rect 209870 200767 209926 200776
rect 302332 200796 302384 200802
rect 209884 200734 209912 200767
rect 302332 200738 302384 200744
rect 209872 200728 209924 200734
rect 209872 200670 209924 200676
rect 204352 200660 204404 200666
rect 204352 200602 204404 200608
rect 204260 200592 204312 200598
rect 201314 200560 201370 200569
rect 200120 200524 200172 200530
rect 201314 200495 201370 200504
rect 201498 200560 201554 200569
rect 201498 200495 201554 200504
rect 201866 200560 201922 200569
rect 204260 200534 204312 200540
rect 201866 200495 201922 200504
rect 200120 200466 200172 200472
rect 198740 200388 198792 200394
rect 198740 200330 198792 200336
rect 197360 200320 197412 200326
rect 197360 200262 197412 200268
rect 196164 200252 196216 200258
rect 196164 200194 196216 200200
rect 201132 200252 201184 200258
rect 201132 200194 201184 200200
rect 178684 200184 178736 200190
rect 201144 200161 201172 200194
rect 201328 200161 201356 200495
rect 201512 200462 201540 200495
rect 201500 200456 201552 200462
rect 201500 200398 201552 200404
rect 201880 200258 201908 200495
rect 220818 200288 220874 200297
rect 201868 200252 201920 200258
rect 220818 200223 220874 200232
rect 201868 200194 201920 200200
rect 220832 200190 220860 200223
rect 220820 200184 220872 200190
rect 178684 200126 178736 200132
rect 201130 200152 201186 200161
rect 201130 200087 201186 200096
rect 201314 200152 201370 200161
rect 220820 200126 220872 200132
rect 201314 200087 201370 200096
rect 318076 13326 318104 256158
rect 318798 220824 318854 220833
rect 318798 220759 318854 220768
rect 318812 220425 318840 220759
rect 318798 220416 318854 220425
rect 318798 220351 318854 220360
rect 318812 203862 318840 220351
rect 318890 218920 318946 218929
rect 318890 218855 318946 218864
rect 318904 218113 318932 218855
rect 318890 218104 318946 218113
rect 318890 218039 318946 218048
rect 318904 204066 318932 218039
rect 319456 217705 319484 261462
rect 319548 260302 319576 341663
rect 319626 340096 319682 340105
rect 319626 340031 319682 340040
rect 319536 260296 319588 260302
rect 319536 260238 319588 260244
rect 319640 260166 319668 340031
rect 319718 338736 319774 338745
rect 319718 338671 319774 338680
rect 319732 260234 319760 338671
rect 319810 337240 319866 337249
rect 319810 337175 319866 337184
rect 319824 261594 319852 337175
rect 319902 336016 319958 336025
rect 319902 335951 319958 335960
rect 319916 262206 319944 335951
rect 319904 262200 319956 262206
rect 319904 262142 319956 262148
rect 319812 261588 319864 261594
rect 319812 261530 319864 261536
rect 319720 260228 319772 260234
rect 319720 260170 319772 260176
rect 319628 260160 319680 260166
rect 319628 260102 319680 260108
rect 319640 221785 319668 260102
rect 319626 221776 319682 221785
rect 319626 221711 319682 221720
rect 319732 220833 319760 260170
rect 319718 220824 319774 220833
rect 319718 220759 319774 220768
rect 319824 218113 319852 261530
rect 319904 223576 319956 223582
rect 319904 223518 319956 223524
rect 319916 223417 319944 223518
rect 319902 223408 319958 223417
rect 319902 223343 319958 223352
rect 319810 218104 319866 218113
rect 319810 218039 319866 218048
rect 319442 217696 319498 217705
rect 319442 217631 319498 217640
rect 318892 204060 318944 204066
rect 318892 204002 318944 204008
rect 318800 203856 318852 203862
rect 318800 203798 318852 203804
rect 320836 44878 320864 397462
rect 320928 385014 320956 500958
rect 321008 408740 321060 408746
rect 321008 408682 321060 408688
rect 320916 385008 320968 385014
rect 320916 384950 320968 384956
rect 320916 358828 320968 358834
rect 320916 358770 320968 358776
rect 320928 290154 320956 358770
rect 321020 306338 321048 408682
rect 321376 407448 321428 407454
rect 321376 407390 321428 407396
rect 321098 406328 321154 406337
rect 321098 406263 321154 406272
rect 321112 325650 321140 406263
rect 321284 405884 321336 405890
rect 321284 405826 321336 405832
rect 321192 394732 321244 394738
rect 321192 394674 321244 394680
rect 321100 325644 321152 325650
rect 321100 325586 321152 325592
rect 321204 321065 321232 394674
rect 321296 336734 321324 405826
rect 321388 371210 321416 407390
rect 322216 401130 322244 572902
rect 323584 572892 323636 572898
rect 323584 572834 323636 572840
rect 322296 553444 322348 553450
rect 322296 553386 322348 553392
rect 322204 401124 322256 401130
rect 322204 401066 322256 401072
rect 322204 396092 322256 396098
rect 322204 396034 322256 396040
rect 321376 371204 321428 371210
rect 321376 371146 321428 371152
rect 321284 336728 321336 336734
rect 321284 336670 321336 336676
rect 321284 334008 321336 334014
rect 321284 333950 321336 333956
rect 321190 321056 321246 321065
rect 321190 320991 321246 321000
rect 321008 306332 321060 306338
rect 321008 306274 321060 306280
rect 321008 294636 321060 294642
rect 321008 294578 321060 294584
rect 320916 290148 320968 290154
rect 320916 290090 320968 290096
rect 320916 288448 320968 288454
rect 320916 288390 320968 288396
rect 320928 270434 320956 288390
rect 321020 284306 321048 294578
rect 321296 292330 321324 333950
rect 321284 292324 321336 292330
rect 321284 292266 321336 292272
rect 322020 289468 322072 289474
rect 322020 289410 322072 289416
rect 321008 284300 321060 284306
rect 321008 284242 321060 284248
rect 322032 281450 322060 289410
rect 322020 281444 322072 281450
rect 322020 281386 322072 281392
rect 320916 270428 320968 270434
rect 320916 270370 320968 270376
rect 320916 256352 320968 256358
rect 320916 256294 320968 256300
rect 320824 44872 320876 44878
rect 320824 44814 320876 44820
rect 318064 13320 318116 13326
rect 318064 13262 318116 13268
rect 124128 10328 124180 10334
rect 124128 10270 124180 10276
rect 122288 4820 122340 4826
rect 122288 4762 122340 4768
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 480 122328 4762
rect 124140 3738 124168 10270
rect 320928 9246 320956 256294
rect 322216 20670 322244 396034
rect 322308 383654 322336 553386
rect 322754 409456 322810 409465
rect 322754 409391 322810 409400
rect 322572 408536 322624 408542
rect 322572 408478 322624 408484
rect 322388 405952 322440 405958
rect 322388 405894 322440 405900
rect 322296 383648 322348 383654
rect 322296 383590 322348 383596
rect 322296 361616 322348 361622
rect 322296 361558 322348 361564
rect 322308 290902 322336 361558
rect 322400 331226 322428 405894
rect 322480 389224 322532 389230
rect 322480 389166 322532 389172
rect 322388 331220 322440 331226
rect 322388 331162 322440 331168
rect 322388 327140 322440 327146
rect 322388 327082 322440 327088
rect 322400 292262 322428 327082
rect 322492 320929 322520 389166
rect 322584 369850 322612 408478
rect 322664 407652 322716 407658
rect 322664 407594 322716 407600
rect 322676 373998 322704 407594
rect 322768 384946 322796 409391
rect 323596 401402 323624 572834
rect 323584 401396 323636 401402
rect 323584 401338 323636 401344
rect 323584 393372 323636 393378
rect 323584 393314 323636 393320
rect 322756 384940 322808 384946
rect 322756 384882 322808 384888
rect 322664 373992 322716 373998
rect 322664 373934 322716 373940
rect 322572 369844 322624 369850
rect 322572 369786 322624 369792
rect 322572 362976 322624 362982
rect 322572 362918 322624 362924
rect 322478 320920 322534 320929
rect 322478 320855 322534 320864
rect 322584 319938 322612 362918
rect 322664 342304 322716 342310
rect 322664 342246 322716 342252
rect 322572 319932 322624 319938
rect 322572 319874 322624 319880
rect 322676 318646 322704 342246
rect 322664 318640 322716 318646
rect 322664 318582 322716 318588
rect 322388 292256 322440 292262
rect 322388 292198 322440 292204
rect 322480 292188 322532 292194
rect 322480 292130 322532 292136
rect 322296 290896 322348 290902
rect 322296 290838 322348 290844
rect 322296 287292 322348 287298
rect 322296 287234 322348 287240
rect 322308 274650 322336 287234
rect 322492 285666 322520 292130
rect 322480 285660 322532 285666
rect 322480 285602 322532 285608
rect 322296 274644 322348 274650
rect 322296 274586 322348 274592
rect 322296 256148 322348 256154
rect 322296 256090 322348 256096
rect 322204 20664 322256 20670
rect 322204 20606 322256 20612
rect 320916 9240 320968 9246
rect 320916 9182 320968 9188
rect 124680 7608 124732 7614
rect 124680 7550 124732 7556
rect 123484 3732 123536 3738
rect 123484 3674 123536 3680
rect 124128 3732 124180 3738
rect 124128 3674 124180 3680
rect 123496 480 123524 3674
rect 124692 480 124720 7550
rect 322308 3058 322336 256090
rect 323596 97986 323624 393314
rect 323688 380798 323716 670686
rect 336096 656940 336148 656946
rect 336096 656882 336148 656888
rect 331864 576156 331916 576162
rect 331864 576098 331916 576104
rect 327724 573164 327776 573170
rect 327724 573106 327776 573112
rect 324964 572824 325016 572830
rect 324964 572766 325016 572772
rect 324044 409012 324096 409018
rect 324044 408954 324096 408960
rect 323860 407992 323912 407998
rect 323860 407934 323912 407940
rect 323768 401668 323820 401674
rect 323768 401610 323820 401616
rect 323676 380792 323728 380798
rect 323676 380734 323728 380740
rect 323676 351960 323728 351966
rect 323676 351902 323728 351908
rect 323688 292398 323716 351902
rect 323676 292392 323728 292398
rect 323676 292334 323728 292340
rect 323780 271794 323808 401610
rect 323872 333266 323900 407934
rect 323952 406564 324004 406570
rect 323952 406506 324004 406512
rect 323964 335306 323992 406506
rect 324056 349110 324084 408954
rect 324976 401334 325004 572766
rect 325332 448588 325384 448594
rect 325332 448530 325384 448536
rect 325148 410100 325200 410106
rect 325148 410042 325200 410048
rect 324964 401328 325016 401334
rect 324964 401270 325016 401276
rect 325056 392012 325108 392018
rect 325056 391954 325108 391960
rect 324964 390584 325016 390590
rect 324964 390526 325016 390532
rect 324044 349104 324096 349110
rect 324044 349046 324096 349052
rect 324044 343664 324096 343670
rect 324044 343606 324096 343612
rect 323952 335300 324004 335306
rect 323952 335242 324004 335248
rect 323860 333260 323912 333266
rect 323860 333202 323912 333208
rect 323952 332648 324004 332654
rect 323952 332590 324004 332596
rect 323964 321298 323992 332590
rect 323952 321292 324004 321298
rect 323952 321234 324004 321240
rect 323860 318504 323912 318510
rect 323860 318446 323912 318452
rect 323872 285598 323900 318446
rect 324056 318170 324084 343606
rect 324044 318164 324096 318170
rect 324044 318106 324096 318112
rect 324320 289400 324372 289406
rect 324320 289342 324372 289348
rect 323860 285592 323912 285598
rect 323860 285534 323912 285540
rect 324332 282878 324360 289342
rect 324976 289105 325004 390526
rect 324962 289096 325018 289105
rect 324962 289031 325018 289040
rect 324320 282872 324372 282878
rect 324320 282814 324372 282820
rect 323768 271788 323820 271794
rect 323768 271730 323820 271736
rect 323676 256080 323728 256086
rect 323676 256022 323728 256028
rect 323584 97980 323636 97986
rect 323584 97922 323636 97928
rect 322296 3052 322348 3058
rect 322296 2994 322348 3000
rect 323688 2990 323716 256022
rect 324964 256012 325016 256018
rect 324964 255954 325016 255960
rect 323676 2984 323728 2990
rect 323676 2926 323728 2932
rect 324976 2922 325004 255954
rect 325068 150414 325096 391954
rect 325160 313274 325188 410042
rect 325238 406464 325294 406473
rect 325238 406399 325294 406408
rect 325252 329798 325280 406399
rect 325344 386374 325372 448530
rect 326344 410168 326396 410174
rect 326344 410110 326396 410116
rect 325424 408128 325476 408134
rect 325424 408070 325476 408076
rect 325332 386368 325384 386374
rect 325332 386310 325384 386316
rect 325332 357468 325384 357474
rect 325332 357410 325384 357416
rect 325240 329792 325292 329798
rect 325240 329734 325292 329740
rect 325148 313268 325200 313274
rect 325148 313210 325200 313216
rect 325344 293486 325372 357410
rect 325436 347070 325464 408070
rect 325516 407312 325568 407318
rect 325516 407254 325568 407260
rect 325528 361554 325556 407254
rect 325516 361548 325568 361554
rect 325516 361490 325568 361496
rect 325424 347064 325476 347070
rect 325424 347006 325476 347012
rect 325516 346452 325568 346458
rect 325516 346394 325568 346400
rect 325332 293480 325384 293486
rect 325332 293422 325384 293428
rect 325148 293412 325200 293418
rect 325148 293354 325200 293360
rect 325160 276010 325188 293354
rect 325528 292058 325556 346394
rect 326356 318646 326384 410110
rect 326528 409080 326580 409086
rect 326528 409022 326580 409028
rect 326436 406632 326488 406638
rect 326436 406574 326488 406580
rect 326448 338094 326476 406574
rect 326540 351898 326568 409022
rect 327736 401198 327764 573106
rect 330576 462392 330628 462398
rect 330576 462334 330628 462340
rect 327908 410236 327960 410242
rect 327908 410178 327960 410184
rect 327816 407720 327868 407726
rect 327816 407662 327868 407668
rect 327724 401192 327776 401198
rect 327724 401134 327776 401140
rect 327724 389292 327776 389298
rect 327724 389234 327776 389240
rect 326620 372632 326672 372638
rect 326620 372574 326672 372580
rect 326528 351892 326580 351898
rect 326528 351834 326580 351840
rect 326436 338088 326488 338094
rect 326436 338030 326488 338036
rect 326528 336796 326580 336802
rect 326528 336738 326580 336744
rect 326540 321434 326568 336738
rect 326528 321428 326580 321434
rect 326528 321370 326580 321376
rect 326632 318782 326660 372574
rect 326620 318776 326672 318782
rect 326620 318718 326672 318724
rect 326344 318640 326396 318646
rect 326344 318582 326396 318588
rect 327736 293962 327764 389234
rect 327828 300830 327856 407662
rect 327920 321570 327948 410178
rect 329196 410032 329248 410038
rect 329196 409974 329248 409980
rect 328276 409760 328328 409766
rect 328276 409702 328328 409708
rect 328000 408332 328052 408338
rect 328000 408274 328052 408280
rect 328012 378146 328040 408274
rect 328184 407380 328236 407386
rect 328184 407322 328236 407328
rect 328092 389360 328144 389366
rect 328092 389302 328144 389308
rect 328000 378140 328052 378146
rect 328000 378082 328052 378088
rect 328000 364404 328052 364410
rect 328000 364346 328052 364352
rect 327908 321564 327960 321570
rect 327908 321506 327960 321512
rect 327908 312588 327960 312594
rect 327908 312530 327960 312536
rect 327816 300824 327868 300830
rect 327816 300766 327868 300772
rect 327724 293956 327776 293962
rect 327724 293898 327776 293904
rect 327816 293548 327868 293554
rect 327816 293490 327868 293496
rect 325516 292052 325568 292058
rect 325516 291994 325568 292000
rect 327724 289672 327776 289678
rect 327724 289614 327776 289620
rect 325148 276004 325200 276010
rect 325148 275946 325200 275952
rect 327736 259350 327764 289614
rect 327828 262954 327856 293490
rect 327920 284238 327948 312530
rect 328012 293282 328040 364346
rect 328104 320793 328132 389302
rect 328196 362914 328224 407322
rect 328288 387802 328316 409702
rect 329104 394800 329156 394806
rect 329104 394742 329156 394748
rect 328276 387796 328328 387802
rect 328276 387738 328328 387744
rect 328184 362908 328236 362914
rect 328184 362850 328236 362856
rect 328184 349172 328236 349178
rect 328184 349114 328236 349120
rect 328090 320784 328146 320793
rect 328090 320719 328146 320728
rect 328196 318238 328224 349114
rect 328184 318232 328236 318238
rect 328184 318174 328236 318180
rect 328000 293276 328052 293282
rect 328000 293218 328052 293224
rect 327908 284232 327960 284238
rect 327908 284174 327960 284180
rect 327816 262948 327868 262954
rect 327816 262890 327868 262896
rect 327724 259344 327776 259350
rect 327724 259286 327776 259292
rect 327724 256556 327776 256562
rect 327724 256498 327776 256504
rect 325056 150408 325108 150414
rect 325056 150350 325108 150356
rect 327736 3262 327764 256498
rect 329116 137290 329144 394742
rect 329208 315994 329236 409974
rect 329564 409896 329616 409902
rect 329564 409838 329616 409844
rect 329288 408808 329340 408814
rect 329288 408750 329340 408756
rect 329300 343534 329328 408750
rect 329378 407688 329434 407697
rect 329378 407623 329434 407632
rect 329392 353258 329420 407623
rect 329472 407516 329524 407522
rect 329472 407458 329524 407464
rect 329484 379506 329512 407458
rect 329576 387734 329604 409838
rect 330484 393440 330536 393446
rect 330484 393382 330536 393388
rect 329564 387728 329616 387734
rect 329564 387670 329616 387676
rect 329472 379500 329524 379506
rect 329472 379442 329524 379448
rect 329472 367124 329524 367130
rect 329472 367066 329524 367072
rect 329380 353252 329432 353258
rect 329380 353194 329432 353200
rect 329288 343528 329340 343534
rect 329288 343470 329340 343476
rect 329380 332716 329432 332722
rect 329380 332658 329432 332664
rect 329288 322992 329340 322998
rect 329288 322934 329340 322940
rect 329196 315988 329248 315994
rect 329196 315930 329248 315936
rect 329300 291922 329328 322934
rect 329392 321026 329420 332658
rect 329484 321230 329512 367066
rect 329564 360256 329616 360262
rect 329564 360198 329616 360204
rect 329472 321224 329524 321230
rect 329472 321166 329524 321172
rect 329380 321020 329432 321026
rect 329380 320962 329432 320968
rect 329576 319802 329604 360198
rect 329564 319796 329616 319802
rect 329564 319738 329616 319744
rect 329288 291916 329340 291922
rect 329288 291858 329340 291864
rect 329196 291848 329248 291854
rect 329196 291790 329248 291796
rect 329208 277302 329236 291790
rect 329196 277296 329248 277302
rect 329196 277238 329248 277244
rect 330496 188358 330524 393382
rect 330588 386102 330616 462334
rect 330942 409320 330998 409329
rect 330942 409255 330998 409264
rect 330760 408876 330812 408882
rect 330760 408818 330812 408824
rect 330666 406192 330722 406201
rect 330666 406127 330722 406136
rect 330576 386096 330628 386102
rect 330576 386038 330628 386044
rect 330576 375420 330628 375426
rect 330576 375362 330628 375368
rect 330588 291786 330616 375362
rect 330680 327078 330708 406127
rect 330772 346390 330800 408818
rect 330852 407788 330904 407794
rect 330852 407730 330904 407736
rect 330864 354142 330892 407730
rect 330956 382158 330984 409255
rect 331876 382226 331904 576098
rect 331956 573096 332008 573102
rect 331956 573038 332008 573044
rect 331968 400722 331996 573038
rect 334716 573028 334768 573034
rect 334716 572970 334768 572976
rect 334624 565888 334676 565894
rect 334624 565830 334676 565836
rect 332048 409964 332100 409970
rect 332048 409906 332100 409912
rect 331956 400716 332008 400722
rect 331956 400658 332008 400664
rect 331956 392080 332008 392086
rect 331956 392022 332008 392028
rect 331864 382220 331916 382226
rect 331864 382162 331916 382168
rect 330944 382152 330996 382158
rect 330944 382094 330996 382100
rect 330852 354136 330904 354142
rect 330852 354078 330904 354084
rect 331864 352028 331916 352034
rect 331864 351970 331916 351976
rect 330852 350600 330904 350606
rect 330852 350542 330904 350548
rect 330760 346384 330812 346390
rect 330760 346326 330812 346332
rect 330760 335368 330812 335374
rect 330760 335310 330812 335316
rect 330668 327072 330720 327078
rect 330668 327014 330720 327020
rect 330772 321094 330800 335310
rect 330760 321088 330812 321094
rect 330760 321030 330812 321036
rect 330864 318714 330892 350542
rect 331128 325712 331180 325718
rect 331128 325654 331180 325660
rect 331140 320958 331168 325654
rect 331128 320952 331180 320958
rect 331128 320894 331180 320900
rect 330852 318708 330904 318714
rect 330852 318650 330904 318656
rect 330668 318436 330720 318442
rect 330668 318378 330720 318384
rect 330576 291780 330628 291786
rect 330576 291722 330628 291728
rect 330680 278662 330708 318378
rect 331876 291106 331904 351970
rect 331864 291100 331916 291106
rect 331864 291042 331916 291048
rect 331864 289332 331916 289338
rect 331864 289274 331916 289280
rect 330668 278656 330720 278662
rect 330668 278598 330720 278604
rect 331876 277370 331904 289274
rect 331864 277364 331916 277370
rect 331864 277306 331916 277312
rect 331864 256488 331916 256494
rect 331864 256430 331916 256436
rect 330484 188352 330536 188358
rect 330484 188294 330536 188300
rect 329104 137284 329156 137290
rect 329104 137226 329156 137232
rect 327724 3256 327776 3262
rect 327724 3198 327776 3204
rect 331876 3194 331904 256430
rect 331968 203794 331996 392022
rect 332060 310486 332088 409906
rect 333244 409828 333296 409834
rect 333244 409770 333296 409776
rect 332416 408468 332468 408474
rect 332416 408410 332468 408416
rect 332232 407924 332284 407930
rect 332232 407866 332284 407872
rect 332140 406428 332192 406434
rect 332140 406370 332192 406376
rect 332152 332586 332180 406370
rect 332244 339454 332272 407866
rect 332324 406768 332376 406774
rect 332324 406710 332376 406716
rect 332336 350538 332364 406710
rect 332428 365702 332456 408410
rect 332416 365696 332468 365702
rect 332416 365638 332468 365644
rect 332416 354748 332468 354754
rect 332416 354690 332468 354696
rect 332324 350532 332376 350538
rect 332324 350474 332376 350480
rect 332232 339448 332284 339454
rect 332232 339390 332284 339396
rect 332324 338156 332376 338162
rect 332324 338098 332376 338104
rect 332140 332580 332192 332586
rect 332140 332522 332192 332528
rect 332140 328500 332192 328506
rect 332140 328442 332192 328448
rect 332048 310480 332100 310486
rect 332048 310422 332100 310428
rect 332048 292120 332100 292126
rect 332048 292062 332100 292068
rect 332060 282810 332088 292062
rect 332152 291990 332180 328442
rect 332336 321162 332364 338098
rect 332324 321156 332376 321162
rect 332324 321098 332376 321104
rect 332428 319666 332456 354690
rect 332416 319660 332468 319666
rect 332416 319602 332468 319608
rect 333256 303618 333284 409770
rect 333334 408232 333390 408241
rect 333334 408167 333390 408176
rect 333348 343602 333376 408167
rect 334636 383586 334664 565830
rect 334728 401470 334756 572970
rect 335268 409488 335320 409494
rect 335268 409430 335320 409436
rect 334900 407856 334952 407862
rect 334900 407798 334952 407804
rect 334806 407280 334862 407289
rect 334806 407215 334862 407224
rect 334716 401464 334768 401470
rect 334716 401406 334768 401412
rect 334716 390652 334768 390658
rect 334716 390594 334768 390600
rect 334624 383580 334676 383586
rect 334624 383522 334676 383528
rect 333428 368552 333480 368558
rect 333428 368494 333480 368500
rect 333336 343596 333388 343602
rect 333336 343538 333388 343544
rect 333336 339516 333388 339522
rect 333336 339458 333388 339464
rect 333348 318578 333376 339458
rect 333440 319870 333468 368494
rect 334624 353320 334676 353326
rect 334624 353262 334676 353268
rect 333428 319864 333480 319870
rect 333428 319806 333480 319812
rect 333336 318572 333388 318578
rect 333336 318514 333388 318520
rect 333244 303612 333296 303618
rect 333244 303554 333296 303560
rect 332140 291984 332192 291990
rect 332140 291926 332192 291932
rect 334636 291038 334664 353262
rect 334624 291032 334676 291038
rect 334624 290974 334676 290980
rect 334624 287904 334676 287910
rect 334624 287846 334676 287852
rect 332048 282804 332100 282810
rect 332048 282746 332100 282752
rect 334636 278730 334664 287846
rect 334624 278724 334676 278730
rect 334624 278666 334676 278672
rect 334624 256420 334676 256426
rect 334624 256362 334676 256368
rect 331956 203788 332008 203794
rect 331956 203730 332008 203736
rect 331864 3188 331916 3194
rect 331864 3130 331916 3136
rect 334636 3126 334664 256362
rect 334728 202774 334756 390594
rect 334820 320142 334848 407215
rect 334912 331158 334940 407798
rect 335082 407552 335138 407561
rect 335082 407487 335138 407496
rect 334992 406700 335044 406706
rect 334992 406642 335044 406648
rect 335004 347342 335032 406642
rect 335096 358766 335124 407487
rect 335176 365764 335228 365770
rect 335176 365706 335228 365712
rect 335084 358760 335136 358766
rect 335084 358702 335136 358708
rect 334992 347336 335044 347342
rect 334992 347278 335044 347284
rect 334992 345092 335044 345098
rect 334992 345034 335044 345040
rect 334900 331152 334952 331158
rect 334900 331094 334952 331100
rect 335004 321366 335032 345034
rect 335084 329860 335136 329866
rect 335084 329802 335136 329808
rect 334992 321360 335044 321366
rect 334992 321302 335044 321308
rect 334808 320136 334860 320142
rect 334808 320078 334860 320084
rect 334808 318368 334860 318374
rect 334808 318310 334860 318316
rect 334820 275942 334848 318310
rect 335096 315314 335124 329802
rect 335188 319734 335216 365706
rect 335280 364342 335308 409430
rect 336002 396264 336058 396273
rect 336002 396199 336058 396208
rect 335268 364336 335320 364342
rect 335268 364278 335320 364284
rect 335176 319728 335228 319734
rect 335176 319670 335228 319676
rect 335084 315308 335136 315314
rect 335084 315250 335136 315256
rect 334808 275936 334860 275942
rect 334808 275878 334860 275884
rect 334716 202768 334768 202774
rect 334716 202710 334768 202716
rect 336016 84862 336044 396199
rect 336108 380905 336136 656882
rect 454040 627224 454092 627230
rect 454040 627166 454092 627172
rect 454052 626618 454080 627166
rect 454040 626612 454092 626618
rect 454040 626554 454092 626560
rect 451280 618928 451332 618934
rect 451280 618870 451332 618876
rect 452200 618928 452252 618934
rect 452200 618870 452252 618876
rect 449900 610632 449952 610638
rect 449900 610574 449952 610580
rect 449912 610026 449940 610574
rect 449900 610020 449952 610026
rect 449900 609962 449952 609968
rect 447140 602404 447192 602410
rect 447140 602346 447192 602352
rect 447152 601730 447180 602346
rect 447140 601724 447192 601730
rect 447140 601666 447192 601672
rect 445024 589348 445076 589354
rect 445024 589290 445076 589296
rect 445036 578202 445064 589290
rect 444380 578196 444432 578202
rect 444380 578138 444432 578144
rect 445024 578196 445076 578202
rect 445024 578138 445076 578144
rect 444392 577658 444420 578138
rect 444380 577652 444432 577658
rect 444380 577594 444432 577600
rect 339408 576224 339460 576230
rect 339408 576166 339460 576172
rect 339420 575482 339448 576166
rect 339408 575476 339460 575482
rect 339408 575418 339460 575424
rect 337568 409624 337620 409630
rect 337568 409566 337620 409572
rect 336556 409556 336608 409562
rect 336556 409498 336608 409504
rect 336280 408060 336332 408066
rect 336280 408002 336332 408008
rect 336188 406496 336240 406502
rect 336188 406438 336240 406444
rect 336094 380896 336150 380905
rect 336094 380831 336150 380840
rect 336094 357096 336150 357105
rect 336094 357031 336150 357040
rect 336108 291174 336136 357031
rect 336200 339833 336228 406438
rect 336292 342718 336320 408002
rect 336370 407416 336426 407425
rect 336370 407351 336426 407360
rect 336384 355201 336412 407351
rect 336462 371240 336518 371249
rect 336462 371175 336518 371184
rect 336370 355192 336426 355201
rect 336370 355127 336426 355136
rect 336370 348120 336426 348129
rect 336370 348055 336426 348064
rect 336280 342712 336332 342718
rect 336280 342654 336332 342660
rect 336278 341728 336334 341737
rect 336278 341663 336334 341672
rect 336186 339824 336242 339833
rect 336186 339759 336242 339768
rect 336186 331528 336242 331537
rect 336186 331463 336242 331472
rect 336200 320890 336228 331463
rect 336188 320884 336240 320890
rect 336188 320826 336240 320832
rect 336188 318300 336240 318306
rect 336188 318242 336240 318248
rect 336096 291168 336148 291174
rect 336096 291110 336148 291116
rect 336200 270473 336228 318242
rect 336292 318102 336320 341663
rect 336384 319462 336412 348055
rect 336476 322250 336504 371175
rect 336568 366761 336596 409498
rect 337476 408944 337528 408950
rect 337476 408886 337528 408892
rect 337384 408672 337436 408678
rect 337384 408614 337436 408620
rect 336924 382220 336976 382226
rect 336924 382162 336976 382168
rect 336936 381585 336964 382162
rect 336922 381576 336978 381585
rect 336922 381511 336978 381520
rect 336924 380724 336976 380730
rect 336924 380666 336976 380672
rect 336936 379681 336964 380666
rect 336922 379672 336978 379681
rect 336922 379607 336978 379616
rect 337290 377632 337346 377641
rect 337290 377567 337346 377576
rect 337304 376786 337332 377567
rect 337292 376780 337344 376786
rect 337292 376722 337344 376728
rect 337106 376408 337162 376417
rect 337106 376343 337162 376352
rect 337120 375426 337148 376343
rect 337108 375420 337160 375426
rect 337108 375362 337160 375368
rect 336922 372600 336978 372609
rect 336922 372535 336978 372544
rect 336936 371278 336964 372535
rect 336924 371272 336976 371278
rect 336924 371214 336976 371220
rect 337292 369844 337344 369850
rect 337292 369786 337344 369792
rect 337304 369345 337332 369786
rect 337290 369336 337346 369345
rect 337290 369271 337346 369280
rect 336554 366752 336610 366761
rect 336554 366687 336610 366696
rect 337290 366072 337346 366081
rect 337290 366007 337346 366016
rect 337304 365770 337332 366007
rect 337292 365764 337344 365770
rect 337292 365706 337344 365712
rect 337106 362264 337162 362273
rect 337106 362199 337162 362208
rect 337120 361622 337148 362199
rect 337108 361616 337160 361622
rect 337108 361558 337160 361564
rect 336924 361548 336976 361554
rect 336924 361490 336976 361496
rect 336936 360369 336964 361490
rect 336922 360360 336978 360369
rect 336922 360295 336978 360304
rect 336924 358760 336976 358766
rect 336924 358702 336976 358708
rect 336936 357785 336964 358702
rect 336922 357776 336978 357785
rect 336922 357711 336978 357720
rect 336922 353288 336978 353297
rect 336922 353223 336978 353232
rect 336936 351966 336964 353223
rect 337290 352064 337346 352073
rect 337290 351999 337292 352008
rect 337344 351999 337346 352008
rect 337292 351970 337344 351976
rect 336924 351960 336976 351966
rect 336924 351902 336976 351908
rect 336924 347064 336976 347070
rect 336924 347006 336976 347012
rect 336740 342712 336792 342718
rect 336740 342654 336792 342660
rect 336752 338609 336780 342654
rect 336936 341057 336964 347006
rect 336922 341048 336978 341057
rect 336922 340983 336978 340992
rect 337290 340504 337346 340513
rect 337290 340439 337346 340448
rect 337304 339522 337332 340439
rect 337292 339516 337344 339522
rect 337292 339458 337344 339464
rect 337290 339144 337346 339153
rect 337290 339079 337346 339088
rect 336738 338600 336794 338609
rect 336738 338535 336794 338544
rect 337304 338162 337332 339079
rect 337292 338156 337344 338162
rect 337292 338098 337344 338104
rect 337106 327584 337162 327593
rect 337106 327519 337162 327528
rect 337120 327146 337148 327519
rect 337108 327140 337160 327146
rect 337108 327082 337160 327088
rect 336464 322244 336516 322250
rect 336464 322186 336516 322192
rect 336924 321564 336976 321570
rect 336924 321506 336976 321512
rect 336936 320521 336964 321506
rect 336922 320512 336978 320521
rect 336922 320447 336978 320456
rect 336372 319456 336424 319462
rect 336372 319398 336424 319404
rect 336922 318608 336978 318617
rect 336922 318543 336978 318552
rect 336280 318096 336332 318102
rect 336280 318038 336332 318044
rect 336936 317490 336964 318543
rect 336924 317484 336976 317490
rect 336924 317426 336976 317432
rect 337108 310480 337160 310486
rect 337108 310422 337160 310428
rect 337120 310321 337148 310422
rect 337106 310312 337162 310321
rect 337106 310247 337162 310256
rect 337108 309120 337160 309126
rect 337108 309062 337160 309068
rect 337120 308961 337148 309062
rect 337106 308952 337162 308961
rect 337106 308887 337162 308896
rect 337396 307737 337424 408614
rect 337488 359145 337516 408886
rect 337580 371929 337608 409566
rect 337658 397624 337714 397633
rect 337658 397559 337714 397568
rect 337672 397526 337700 397559
rect 337660 397520 337712 397526
rect 337660 397462 337712 397468
rect 337658 396944 337714 396953
rect 337658 396879 337714 396888
rect 337672 396098 337700 396879
rect 337660 396092 337712 396098
rect 337660 396034 337712 396040
rect 337750 395720 337806 395729
rect 337750 395655 337806 395664
rect 337658 395040 337714 395049
rect 337658 394975 337714 394984
rect 337672 394806 337700 394975
rect 337660 394800 337712 394806
rect 337660 394742 337712 394748
rect 337764 394738 337792 395655
rect 337752 394732 337804 394738
rect 337752 394674 337804 394680
rect 337750 394360 337806 394369
rect 337750 394295 337806 394304
rect 337658 393680 337714 393689
rect 337658 393615 337714 393624
rect 337672 393446 337700 393615
rect 337660 393440 337712 393446
rect 337660 393382 337712 393388
rect 337764 393378 337792 394295
rect 337752 393372 337804 393378
rect 337752 393314 337804 393320
rect 337750 393136 337806 393145
rect 337750 393071 337806 393080
rect 337658 392456 337714 392465
rect 337658 392391 337714 392400
rect 337672 392086 337700 392391
rect 337660 392080 337712 392086
rect 337660 392022 337712 392028
rect 337764 392018 337792 393071
rect 337752 392012 337804 392018
rect 337752 391954 337804 391960
rect 337658 391776 337714 391785
rect 337658 391711 337714 391720
rect 337672 390658 337700 391711
rect 337750 391232 337806 391241
rect 337750 391167 337806 391176
rect 337660 390652 337712 390658
rect 337660 390594 337712 390600
rect 337764 390590 337792 391167
rect 337752 390584 337804 390590
rect 337658 390552 337714 390561
rect 337752 390526 337804 390532
rect 337658 390487 337714 390496
rect 337672 389366 337700 390487
rect 337750 389872 337806 389881
rect 337750 389807 337806 389816
rect 337660 389360 337712 389366
rect 337660 389302 337712 389308
rect 337764 389298 337792 389807
rect 337752 389292 337804 389298
rect 337752 389234 337804 389240
rect 337660 389224 337712 389230
rect 337658 389192 337660 389201
rect 337712 389192 337714 389201
rect 337658 389127 337714 389136
rect 337844 389156 337896 389162
rect 337844 389098 337896 389104
rect 337752 389088 337804 389094
rect 337752 389030 337804 389036
rect 337764 388657 337792 389030
rect 337750 388648 337806 388657
rect 337750 388583 337806 388592
rect 337856 387977 337884 389098
rect 337842 387968 337898 387977
rect 337842 387903 337898 387912
rect 337660 387796 337712 387802
rect 337660 387738 337712 387744
rect 337672 387297 337700 387738
rect 337752 387728 337804 387734
rect 337752 387670 337804 387676
rect 337658 387288 337714 387297
rect 337658 387223 337714 387232
rect 337764 386753 337792 387670
rect 337750 386744 337806 386753
rect 337750 386679 337806 386688
rect 337660 386368 337712 386374
rect 337660 386310 337712 386316
rect 337672 386073 337700 386310
rect 337752 386096 337804 386102
rect 337658 386064 337714 386073
rect 337752 386038 337804 386044
rect 337658 385999 337714 386008
rect 337764 385393 337792 386038
rect 337750 385384 337806 385393
rect 337750 385319 337806 385328
rect 337660 385008 337712 385014
rect 337660 384950 337712 384956
rect 337672 384713 337700 384950
rect 337752 384940 337804 384946
rect 337752 384882 337804 384888
rect 337658 384704 337714 384713
rect 337658 384639 337714 384648
rect 337764 384169 337792 384882
rect 337750 384160 337806 384169
rect 337750 384095 337806 384104
rect 337660 383648 337712 383654
rect 337660 383590 337712 383596
rect 337672 383489 337700 383590
rect 337752 383580 337804 383586
rect 337752 383522 337804 383528
rect 337658 383480 337714 383489
rect 337658 383415 337714 383424
rect 337764 382809 337792 383522
rect 337750 382800 337806 382809
rect 337750 382735 337806 382744
rect 337660 382152 337712 382158
rect 337658 382120 337660 382129
rect 337712 382120 337714 382129
rect 337658 382055 337714 382064
rect 337752 380792 337804 380798
rect 337752 380734 337804 380740
rect 337764 380225 337792 380734
rect 337750 380216 337806 380225
rect 337750 380151 337806 380160
rect 337752 379500 337804 379506
rect 337752 379442 337804 379448
rect 337658 378992 337714 379001
rect 337658 378927 337714 378936
rect 337672 378214 337700 378927
rect 337764 378321 337792 379442
rect 337750 378312 337806 378321
rect 337750 378247 337806 378256
rect 337660 378208 337712 378214
rect 337660 378150 337712 378156
rect 337752 378140 337804 378146
rect 337752 378082 337804 378088
rect 337764 377097 337792 378082
rect 337750 377088 337806 377097
rect 337750 377023 337806 377032
rect 337660 376712 337712 376718
rect 337660 376654 337712 376660
rect 337672 375737 337700 376654
rect 337658 375728 337714 375737
rect 337658 375663 337714 375672
rect 337660 375352 337712 375358
rect 337660 375294 337712 375300
rect 337672 374513 337700 375294
rect 337750 375184 337806 375193
rect 337750 375119 337806 375128
rect 337658 374504 337714 374513
rect 337658 374439 337714 374448
rect 337764 374066 337792 375119
rect 337752 374060 337804 374066
rect 337752 374002 337804 374008
rect 337660 373992 337712 373998
rect 337660 373934 337712 373940
rect 337672 373153 337700 373934
rect 337750 373824 337806 373833
rect 337750 373759 337806 373768
rect 337658 373144 337714 373153
rect 337658 373079 337714 373088
rect 337764 372638 337792 373759
rect 337752 372632 337804 372638
rect 337752 372574 337804 372580
rect 337566 371920 337622 371929
rect 337566 371855 337622 371864
rect 337568 371816 337620 371822
rect 337568 371758 337620 371764
rect 337580 361593 337608 371758
rect 337660 371204 337712 371210
rect 337660 371146 337712 371152
rect 337672 370705 337700 371146
rect 337658 370696 337714 370705
rect 337658 370631 337714 370640
rect 337658 370016 337714 370025
rect 337658 369951 337714 369960
rect 337672 369918 337700 369951
rect 337660 369912 337712 369918
rect 337660 369854 337712 369860
rect 337658 368656 337714 368665
rect 337658 368591 337714 368600
rect 337672 368558 337700 368591
rect 337660 368552 337712 368558
rect 337660 368494 337712 368500
rect 337752 368484 337804 368490
rect 337752 368426 337804 368432
rect 337764 368121 337792 368426
rect 337750 368112 337806 368121
rect 337750 368047 337806 368056
rect 337750 367432 337806 367441
rect 337750 367367 337806 367376
rect 337764 367130 337792 367367
rect 337752 367124 337804 367130
rect 337752 367066 337804 367072
rect 337660 365696 337712 365702
rect 337660 365638 337712 365644
rect 337672 365537 337700 365638
rect 337658 365528 337714 365537
rect 337658 365463 337714 365472
rect 337750 364848 337806 364857
rect 337750 364783 337806 364792
rect 337764 364410 337792 364783
rect 337752 364404 337804 364410
rect 337752 364346 337804 364352
rect 337660 364336 337712 364342
rect 337660 364278 337712 364284
rect 337672 364177 337700 364278
rect 337658 364168 337714 364177
rect 337658 364103 337714 364112
rect 337750 363624 337806 363633
rect 337750 363559 337806 363568
rect 337764 362982 337792 363559
rect 337752 362976 337804 362982
rect 337658 362944 337714 362953
rect 337752 362918 337804 362924
rect 337658 362879 337660 362888
rect 337712 362879 337714 362888
rect 337660 362850 337712 362856
rect 337566 361584 337622 361593
rect 337566 361519 337622 361528
rect 337658 361040 337714 361049
rect 337658 360975 337714 360984
rect 337672 360262 337700 360975
rect 337660 360256 337712 360262
rect 337660 360198 337712 360204
rect 337658 359680 337714 359689
rect 337658 359615 337714 359624
rect 337568 359508 337620 359514
rect 337568 359450 337620 359456
rect 337474 359136 337530 359145
rect 337474 359071 337530 359080
rect 337476 354136 337528 354142
rect 337476 354078 337528 354084
rect 337488 353818 337516 354078
rect 337580 353977 337608 359450
rect 337672 358834 337700 359615
rect 337660 358828 337712 358834
rect 337660 358770 337712 358776
rect 337750 358456 337806 358465
rect 337750 358391 337806 358400
rect 337764 357474 337792 358391
rect 337752 357468 337804 357474
rect 337752 357410 337804 357416
rect 337660 357400 337712 357406
rect 337660 357342 337712 357348
rect 337672 356561 337700 357342
rect 337658 356552 337714 356561
rect 337658 356487 337714 356496
rect 337658 355872 337714 355881
rect 337658 355807 337714 355816
rect 337672 354754 337700 355807
rect 337660 354748 337712 354754
rect 337660 354690 337712 354696
rect 337750 354648 337806 354657
rect 337750 354583 337806 354592
rect 337566 353968 337622 353977
rect 337566 353903 337622 353912
rect 337488 353790 337608 353818
rect 337474 346896 337530 346905
rect 337474 346831 337530 346840
rect 337488 346458 337516 346831
rect 337476 346452 337528 346458
rect 337476 346394 337528 346400
rect 337580 345014 337608 353790
rect 337764 353326 337792 354583
rect 337752 353320 337804 353326
rect 337752 353262 337804 353268
rect 337660 353252 337712 353258
rect 337660 353194 337712 353200
rect 337672 352617 337700 353194
rect 337658 352608 337714 352617
rect 337658 352543 337714 352552
rect 337660 351892 337712 351898
rect 337660 351834 337712 351840
rect 337672 351393 337700 351834
rect 337658 351384 337714 351393
rect 337658 351319 337714 351328
rect 337658 350704 337714 350713
rect 337658 350639 337714 350648
rect 337672 350606 337700 350639
rect 337660 350600 337712 350606
rect 337660 350542 337712 350548
rect 337752 350532 337804 350538
rect 337752 350474 337804 350480
rect 337764 350033 337792 350474
rect 337750 350024 337806 350033
rect 337750 349959 337806 349968
rect 337658 349480 337714 349489
rect 337658 349415 337714 349424
rect 337672 349178 337700 349415
rect 337660 349172 337712 349178
rect 337660 349114 337712 349120
rect 337752 349104 337804 349110
rect 337752 349046 337804 349052
rect 337764 348809 337792 349046
rect 337750 348800 337806 348809
rect 337750 348735 337806 348744
rect 337658 347576 337714 347585
rect 337658 347511 337714 347520
rect 337672 347342 337700 347511
rect 337660 347336 337712 347342
rect 337660 347278 337712 347284
rect 337660 346384 337712 346390
rect 337660 346326 337712 346332
rect 337672 346225 337700 346326
rect 337658 346216 337714 346225
rect 337658 346151 337714 346160
rect 337658 345536 337714 345545
rect 337658 345471 337714 345480
rect 337672 345098 337700 345471
rect 337660 345092 337712 345098
rect 337660 345034 337712 345040
rect 337488 344986 337608 345014
rect 337752 345024 337804 345030
rect 337750 344992 337752 345001
rect 337804 344992 337806 345001
rect 337488 323105 337516 344986
rect 337750 344927 337806 344936
rect 337658 344312 337714 344321
rect 337658 344247 337714 344256
rect 337672 343670 337700 344247
rect 337660 343664 337712 343670
rect 337660 343606 337712 343612
rect 337750 343632 337806 343641
rect 337568 343596 337620 343602
rect 337750 343567 337806 343576
rect 337568 343538 337620 343544
rect 337580 342417 337608 343538
rect 337764 343534 337792 343567
rect 337752 343528 337804 343534
rect 337752 343470 337804 343476
rect 337658 343088 337714 343097
rect 337658 343023 337714 343032
rect 337566 342408 337622 342417
rect 337566 342343 337622 342352
rect 337672 342310 337700 343023
rect 337660 342304 337712 342310
rect 337660 342246 337712 342252
rect 337568 339448 337620 339454
rect 337568 339390 337620 339396
rect 337580 335866 337608 339390
rect 337660 338088 337712 338094
rect 337660 338030 337712 338036
rect 337672 337249 337700 338030
rect 337750 337920 337806 337929
rect 337750 337855 337806 337864
rect 337658 337240 337714 337249
rect 337658 337175 337714 337184
rect 337764 336802 337792 337855
rect 337752 336796 337804 336802
rect 337752 336738 337804 336744
rect 337660 336728 337712 336734
rect 337660 336670 337712 336676
rect 337672 336025 337700 336670
rect 337842 336560 337898 336569
rect 337842 336495 337898 336504
rect 337658 336016 337714 336025
rect 337658 335951 337714 335960
rect 337580 335838 337700 335866
rect 337566 335336 337622 335345
rect 337566 335271 337622 335280
rect 337580 334014 337608 335271
rect 337672 334370 337700 335838
rect 337856 335374 337884 336495
rect 337844 335368 337896 335374
rect 337844 335310 337896 335316
rect 337752 335300 337804 335306
rect 337752 335242 337804 335248
rect 337764 334665 337792 335242
rect 337750 334656 337806 334665
rect 337750 334591 337806 334600
rect 337672 334342 337792 334370
rect 337568 334008 337620 334014
rect 337568 333950 337620 333956
rect 337658 333976 337714 333985
rect 337658 333911 337714 333920
rect 337672 332722 337700 333911
rect 337764 333441 337792 334342
rect 337750 333432 337806 333441
rect 337750 333367 337806 333376
rect 337844 333260 337896 333266
rect 337844 333202 337896 333208
rect 337750 332752 337806 332761
rect 337660 332716 337712 332722
rect 337750 332687 337806 332696
rect 337660 332658 337712 332664
rect 337764 332654 337792 332687
rect 337752 332648 337804 332654
rect 337752 332590 337804 332596
rect 337660 332580 337712 332586
rect 337660 332522 337712 332528
rect 337672 332081 337700 332522
rect 337658 332072 337714 332081
rect 337658 332007 337714 332016
rect 337660 331220 337712 331226
rect 337660 331162 337712 331168
rect 337568 331152 337620 331158
rect 337568 331094 337620 331100
rect 337580 328273 337608 331094
rect 337672 330857 337700 331162
rect 337658 330848 337714 330857
rect 337658 330783 337714 330792
rect 337750 330168 337806 330177
rect 337750 330103 337806 330112
rect 337764 329866 337792 330103
rect 337752 329860 337804 329866
rect 337752 329802 337804 329808
rect 337660 329792 337712 329798
rect 337660 329734 337712 329740
rect 337672 329497 337700 329734
rect 337658 329488 337714 329497
rect 337658 329423 337714 329432
rect 337658 328944 337714 328953
rect 337658 328879 337714 328888
rect 337672 328506 337700 328879
rect 337660 328500 337712 328506
rect 337660 328442 337712 328448
rect 337566 328264 337622 328273
rect 337566 328199 337622 328208
rect 337856 328114 337884 333202
rect 337580 328086 337884 328114
rect 337580 325689 337608 328086
rect 337660 327072 337712 327078
rect 337658 327040 337660 327049
rect 337712 327040 337714 327049
rect 337658 326975 337714 326984
rect 337658 326360 337714 326369
rect 337658 326295 337714 326304
rect 337672 325718 337700 326295
rect 337660 325712 337712 325718
rect 337566 325680 337622 325689
rect 337660 325654 337712 325660
rect 337566 325615 337622 325624
rect 337752 325644 337804 325650
rect 337752 325586 337804 325592
rect 337658 325000 337714 325009
rect 337658 324935 337714 324944
rect 337672 324358 337700 324935
rect 337764 324465 337792 325586
rect 337750 324456 337806 324465
rect 337750 324391 337806 324400
rect 337660 324352 337712 324358
rect 337660 324294 337712 324300
rect 337658 323776 337714 323785
rect 337658 323711 337714 323720
rect 337474 323096 337530 323105
rect 337474 323031 337530 323040
rect 337672 322998 337700 323711
rect 337660 322992 337712 322998
rect 337660 322934 337712 322940
rect 337750 322552 337806 322561
rect 337750 322487 337806 322496
rect 337660 322448 337712 322454
rect 337660 322390 337712 322396
rect 337672 321881 337700 322390
rect 337658 321872 337714 321881
rect 337658 321807 337714 321816
rect 337764 321638 337792 322487
rect 337752 321632 337804 321638
rect 337752 321574 337804 321580
rect 337660 321496 337712 321502
rect 337660 321438 337712 321444
rect 337672 321201 337700 321438
rect 337658 321192 337714 321201
rect 337658 321127 337714 321136
rect 337660 320136 337712 320142
rect 337660 320078 337712 320084
rect 337672 319297 337700 320078
rect 337750 319968 337806 319977
rect 337750 319903 337806 319912
rect 337658 319288 337714 319297
rect 337658 319223 337714 319232
rect 337764 318850 337792 319903
rect 337752 318844 337804 318850
rect 337752 318786 337804 318792
rect 337660 318640 337712 318646
rect 337660 318582 337712 318588
rect 337672 317937 337700 318582
rect 337658 317928 337714 317937
rect 337658 317863 337714 317872
rect 337660 317416 337712 317422
rect 337566 317384 337622 317393
rect 337660 317358 337712 317364
rect 337566 317319 337622 317328
rect 337580 316062 337608 317319
rect 337672 316713 337700 317358
rect 337658 316704 337714 316713
rect 337658 316639 337714 316648
rect 337568 316056 337620 316062
rect 337568 315998 337620 316004
rect 337750 316024 337806 316033
rect 337660 315988 337712 315994
rect 337750 315959 337806 315968
rect 337660 315930 337712 315936
rect 337672 315489 337700 315930
rect 337658 315480 337714 315489
rect 337658 315415 337714 315424
rect 337658 314800 337714 314809
rect 337658 314735 337660 314744
rect 337712 314735 337714 314744
rect 337660 314706 337712 314712
rect 337764 314702 337792 315959
rect 337752 314696 337804 314702
rect 337752 314638 337804 314644
rect 337660 314628 337712 314634
rect 337660 314570 337712 314576
rect 337672 314129 337700 314570
rect 337658 314120 337714 314129
rect 337658 314055 337714 314064
rect 337658 313440 337714 313449
rect 337658 313375 337714 313384
rect 337672 313342 337700 313375
rect 337660 313336 337712 313342
rect 337660 313278 337712 313284
rect 337752 313268 337804 313274
rect 337752 313210 337804 313216
rect 337764 312905 337792 313210
rect 337750 312896 337806 312905
rect 337750 312831 337806 312840
rect 337750 312216 337806 312225
rect 337750 312151 337806 312160
rect 337764 311914 337792 312151
rect 337752 311908 337804 311914
rect 337752 311850 337804 311856
rect 337660 311840 337712 311846
rect 337660 311782 337712 311788
rect 337672 311545 337700 311782
rect 337658 311536 337714 311545
rect 337658 311471 337714 311480
rect 337658 310992 337714 311001
rect 337658 310927 337714 310936
rect 337672 310554 337700 310927
rect 337660 310548 337712 310554
rect 337660 310490 337712 310496
rect 337658 309632 337714 309641
rect 337658 309567 337714 309576
rect 337672 309194 337700 309567
rect 337660 309188 337712 309194
rect 337660 309130 337712 309136
rect 337658 308408 337714 308417
rect 337658 308343 337714 308352
rect 337672 307834 337700 308343
rect 337660 307828 337712 307834
rect 337660 307770 337712 307776
rect 337752 307760 337804 307766
rect 337382 307728 337438 307737
rect 337752 307702 337804 307708
rect 337382 307663 337438 307672
rect 337658 307048 337714 307057
rect 337658 306983 337714 306992
rect 337672 306406 337700 306983
rect 337764 306513 337792 307702
rect 337750 306504 337806 306513
rect 337750 306439 337806 306448
rect 337660 306400 337712 306406
rect 337660 306342 337712 306348
rect 337752 306332 337804 306338
rect 337752 306274 337804 306280
rect 337658 305824 337714 305833
rect 337658 305759 337714 305768
rect 337672 305046 337700 305759
rect 337764 305153 337792 306274
rect 337750 305144 337806 305153
rect 337750 305079 337806 305088
rect 337660 305040 337712 305046
rect 337660 304982 337712 304988
rect 337752 304972 337804 304978
rect 337752 304914 337804 304920
rect 337658 304464 337714 304473
rect 337658 304399 337714 304408
rect 337672 303686 337700 304399
rect 337764 303929 337792 304914
rect 337750 303920 337806 303929
rect 337750 303855 337806 303864
rect 337660 303680 337712 303686
rect 337660 303622 337712 303628
rect 336924 303612 336976 303618
rect 336924 303554 336976 303560
rect 336936 302569 336964 303554
rect 337658 303240 337714 303249
rect 337658 303175 337714 303184
rect 336922 302560 336978 302569
rect 336922 302495 336978 302504
rect 337672 302258 337700 303175
rect 337660 302252 337712 302258
rect 337660 302194 337712 302200
rect 337476 302184 337528 302190
rect 337476 302126 337528 302132
rect 337488 301345 337516 302126
rect 337658 301880 337714 301889
rect 337658 301815 337714 301824
rect 337474 301336 337530 301345
rect 337474 301271 337530 301280
rect 337672 300898 337700 301815
rect 337660 300892 337712 300898
rect 337660 300834 337712 300840
rect 337384 300824 337436 300830
rect 337384 300766 337436 300772
rect 337396 299985 337424 300766
rect 337658 300656 337714 300665
rect 337658 300591 337714 300600
rect 337382 299976 337438 299985
rect 337382 299911 337438 299920
rect 337672 299538 337700 300591
rect 337660 299532 337712 299538
rect 337660 299474 337712 299480
rect 337292 299464 337344 299470
rect 337106 299432 337162 299441
rect 337292 299406 337344 299412
rect 337106 299367 337162 299376
rect 337120 298178 337148 299367
rect 337304 298761 337332 299406
rect 337290 298752 337346 298761
rect 337290 298687 337346 298696
rect 337108 298172 337160 298178
rect 337108 298114 337160 298120
rect 336924 298104 336976 298110
rect 336924 298046 336976 298052
rect 337750 298072 337806 298081
rect 336936 296857 336964 298046
rect 337660 298036 337712 298042
rect 337750 298007 337806 298016
rect 337660 297978 337712 297984
rect 337672 297401 337700 297978
rect 337658 297392 337714 297401
rect 337658 297327 337714 297336
rect 336922 296848 336978 296857
rect 336922 296783 336978 296792
rect 337764 296750 337792 298007
rect 337752 296744 337804 296750
rect 337752 296686 337804 296692
rect 337108 296676 337160 296682
rect 337108 296618 337160 296624
rect 337120 295497 337148 296618
rect 337660 296608 337712 296614
rect 337660 296550 337712 296556
rect 337672 296177 337700 296550
rect 337658 296168 337714 296177
rect 337658 296103 337714 296112
rect 337106 295488 337162 295497
rect 337106 295423 337162 295432
rect 337660 295316 337712 295322
rect 337660 295258 337712 295264
rect 336922 294944 336978 294953
rect 336922 294879 336978 294888
rect 336936 294030 336964 294879
rect 337672 294273 337700 295258
rect 337658 294264 337714 294273
rect 337658 294199 337714 294208
rect 336924 294024 336976 294030
rect 336924 293966 336976 293972
rect 337752 293888 337804 293894
rect 337752 293830 337804 293836
rect 337660 293820 337712 293826
rect 337660 293762 337712 293768
rect 337672 293593 337700 293762
rect 337658 293584 337714 293593
rect 337658 293519 337714 293528
rect 336280 293344 336332 293350
rect 336280 293286 336332 293292
rect 336292 280809 336320 293286
rect 337764 292913 337792 293830
rect 337750 292904 337806 292913
rect 337750 292839 337806 292848
rect 337660 292528 337712 292534
rect 337660 292470 337712 292476
rect 337672 292369 337700 292470
rect 337752 292460 337804 292466
rect 337752 292402 337804 292408
rect 337658 292360 337714 292369
rect 337658 292295 337714 292304
rect 337764 291689 337792 292402
rect 337750 291680 337806 291689
rect 337750 291615 337806 291624
rect 337474 291000 337530 291009
rect 337108 290964 337160 290970
rect 337474 290935 337530 290944
rect 337108 290906 337160 290912
rect 337120 290465 337148 290906
rect 337106 290456 337162 290465
rect 337106 290391 337162 290400
rect 337488 290358 337516 290935
rect 337476 290352 337528 290358
rect 337476 290294 337528 290300
rect 337752 289808 337804 289814
rect 337658 289776 337714 289785
rect 337752 289750 337804 289756
rect 337658 289711 337660 289720
rect 337712 289711 337714 289720
rect 337660 289682 337712 289688
rect 337476 289264 337528 289270
rect 337476 289206 337528 289212
rect 336740 289196 336792 289202
rect 336740 289138 336792 289144
rect 336752 287638 336780 289138
rect 337384 288856 337436 288862
rect 337384 288798 337436 288804
rect 336832 288516 336884 288522
rect 336832 288458 336884 288464
rect 336740 287632 336792 287638
rect 336740 287574 336792 287580
rect 336844 287042 336872 288458
rect 336924 288380 336976 288386
rect 336924 288322 336976 288328
rect 336936 287201 336964 288322
rect 337200 288040 337252 288046
rect 337200 287982 337252 287988
rect 337108 287836 337160 287842
rect 337108 287778 337160 287784
rect 337016 287768 337068 287774
rect 337016 287710 337068 287716
rect 336922 287192 336978 287201
rect 336922 287127 336978 287136
rect 337028 287054 337056 287710
rect 336660 287014 336872 287042
rect 336936 287026 337056 287054
rect 336660 285190 336688 287014
rect 336740 286952 336792 286958
rect 336740 286894 336792 286900
rect 336752 286521 336780 286894
rect 336832 286884 336884 286890
rect 336832 286826 336884 286832
rect 336738 286512 336794 286521
rect 336738 286447 336794 286456
rect 336740 285728 336792 285734
rect 336740 285670 336792 285676
rect 336648 285184 336700 285190
rect 336648 285126 336700 285132
rect 336278 280800 336334 280809
rect 336278 280735 336334 280744
rect 336752 279449 336780 285670
rect 336844 280129 336872 286826
rect 336830 280120 336886 280129
rect 336830 280055 336886 280064
rect 336738 279440 336794 279449
rect 336738 279375 336794 279384
rect 336936 277394 336964 287026
rect 337120 286890 337148 287778
rect 337212 287026 337240 287982
rect 337292 287972 337344 287978
rect 337292 287914 337344 287920
rect 337200 287020 337252 287026
rect 337200 286962 337252 286968
rect 337108 286884 337160 286890
rect 337108 286826 337160 286832
rect 337200 286884 337252 286890
rect 337200 286826 337252 286832
rect 337106 286784 337162 286793
rect 337106 286719 337162 286728
rect 337016 285796 337068 285802
rect 337016 285738 337068 285744
rect 337028 277545 337056 285738
rect 337120 277642 337148 286719
rect 337212 277642 337240 286826
rect 337304 285734 337332 287914
rect 337292 285728 337344 285734
rect 337292 285670 337344 285676
rect 337292 285592 337344 285598
rect 337292 285534 337344 285540
rect 337304 285297 337332 285534
rect 337290 285288 337346 285297
rect 337290 285223 337346 285232
rect 337292 285184 337344 285190
rect 337292 285126 337344 285132
rect 337304 282402 337332 285126
rect 337292 282396 337344 282402
rect 337292 282338 337344 282344
rect 337396 282282 337424 288798
rect 337488 286929 337516 289206
rect 337764 289105 337792 289750
rect 338764 289128 338816 289134
rect 337750 289096 337806 289105
rect 338764 289070 338816 289076
rect 337750 289031 337806 289040
rect 337568 288924 337620 288930
rect 337568 288866 337620 288872
rect 337580 288130 337608 288866
rect 338028 288720 338080 288726
rect 338028 288662 338080 288668
rect 337936 288652 337988 288658
rect 337936 288594 337988 288600
rect 337844 288584 337896 288590
rect 337844 288526 337896 288532
rect 337658 288416 337714 288425
rect 337658 288351 337714 288360
rect 337672 288318 337700 288351
rect 337660 288312 337712 288318
rect 337660 288254 337712 288260
rect 337752 288244 337804 288250
rect 337752 288186 337804 288192
rect 337580 288102 337700 288130
rect 337672 287722 337700 288102
rect 337764 287881 337792 288186
rect 337750 287872 337806 287881
rect 337750 287807 337806 287816
rect 337568 287700 337620 287706
rect 337672 287694 337792 287722
rect 337568 287642 337620 287648
rect 337474 286920 337530 286929
rect 337474 286855 337530 286864
rect 337476 286816 337528 286822
rect 337476 286758 337528 286764
rect 337488 285841 337516 286758
rect 337474 285832 337530 285841
rect 337474 285767 337530 285776
rect 337476 284368 337528 284374
rect 337476 284310 337528 284316
rect 337304 282254 337424 282282
rect 337108 277636 337160 277642
rect 337108 277578 337160 277584
rect 337200 277636 337252 277642
rect 337200 277578 337252 277584
rect 337014 277536 337070 277545
rect 337014 277471 337070 277480
rect 337198 277536 337254 277545
rect 337198 277471 337254 277480
rect 337108 277432 337160 277438
rect 336844 277366 336964 277394
rect 337014 277400 337070 277409
rect 336186 270464 336242 270473
rect 336186 270399 336242 270408
rect 336844 264081 336872 277366
rect 337108 277374 337160 277380
rect 337014 277335 337070 277344
rect 337028 269249 337056 277335
rect 337120 274417 337148 277374
rect 337106 274408 337162 274417
rect 337106 274343 337162 274352
rect 337212 273057 337240 277471
rect 337304 277409 337332 282254
rect 337384 282192 337436 282198
rect 337384 282134 337436 282140
rect 337396 277982 337424 282134
rect 337384 277976 337436 277982
rect 337384 277918 337436 277924
rect 337290 277400 337346 277409
rect 337290 277335 337346 277344
rect 337384 277364 337436 277370
rect 337384 277306 337436 277312
rect 337290 277264 337346 277273
rect 337290 277199 337346 277208
rect 337198 273048 337254 273057
rect 337198 272983 337254 272992
rect 337106 271824 337162 271833
rect 337106 271759 337108 271768
rect 337160 271759 337162 271768
rect 337108 271730 337160 271736
rect 337014 269240 337070 269249
rect 337014 269175 337070 269184
rect 337304 268569 337332 277199
rect 337396 276321 337424 277306
rect 337382 276312 337438 276321
rect 337382 276247 337438 276256
rect 337384 275936 337436 275942
rect 337384 275878 337436 275884
rect 337396 274961 337424 275878
rect 337382 274952 337438 274961
rect 337382 274887 337438 274896
rect 337290 268560 337346 268569
rect 337290 268495 337346 268504
rect 337488 265305 337516 284310
rect 337474 265296 337530 265305
rect 337474 265231 337530 265240
rect 337580 264761 337608 287642
rect 337660 287632 337712 287638
rect 337660 287574 337712 287580
rect 337672 285802 337700 287574
rect 337660 285796 337712 285802
rect 337660 285738 337712 285744
rect 337660 285660 337712 285666
rect 337660 285602 337712 285608
rect 337672 284617 337700 285602
rect 337658 284608 337714 284617
rect 337658 284543 337714 284552
rect 337764 284374 337792 287694
rect 337752 284368 337804 284374
rect 337752 284310 337804 284316
rect 337660 284300 337712 284306
rect 337660 284242 337712 284248
rect 337672 283937 337700 284242
rect 337752 284232 337804 284238
rect 337752 284174 337804 284180
rect 337658 283928 337714 283937
rect 337658 283863 337714 283872
rect 337764 283393 337792 284174
rect 337750 283384 337806 283393
rect 337750 283319 337806 283328
rect 337660 282872 337712 282878
rect 337660 282814 337712 282820
rect 337672 282713 337700 282814
rect 337752 282804 337804 282810
rect 337752 282746 337804 282752
rect 337658 282704 337714 282713
rect 337658 282639 337714 282648
rect 337660 282600 337712 282606
rect 337660 282542 337712 282548
rect 337672 281874 337700 282542
rect 337764 282033 337792 282746
rect 337750 282024 337806 282033
rect 337750 281959 337806 281968
rect 337672 281846 337792 281874
rect 337660 281444 337712 281450
rect 337660 281386 337712 281392
rect 337672 281353 337700 281386
rect 337658 281344 337714 281353
rect 337658 281279 337714 281288
rect 337764 278905 337792 281846
rect 337750 278896 337806 278905
rect 337750 278831 337806 278840
rect 337660 278724 337712 278730
rect 337660 278666 337712 278672
rect 337672 278225 337700 278666
rect 337752 278656 337804 278662
rect 337752 278598 337804 278604
rect 337658 278216 337714 278225
rect 337658 278151 337714 278160
rect 337660 278112 337712 278118
rect 337660 278054 337712 278060
rect 337672 265985 337700 278054
rect 337764 277545 337792 278598
rect 337750 277536 337806 277545
rect 337750 277471 337806 277480
rect 337752 277432 337804 277438
rect 337856 277409 337884 288526
rect 337948 287298 337976 288594
rect 338040 287298 338068 288662
rect 337936 287292 337988 287298
rect 337936 287234 337988 287240
rect 338028 287292 338080 287298
rect 338028 287234 338080 287240
rect 337936 287088 337988 287094
rect 337936 287030 337988 287036
rect 338028 287088 338080 287094
rect 338080 287036 338160 287042
rect 338028 287030 338160 287036
rect 337948 286906 337976 287030
rect 338040 287014 338160 287030
rect 337948 286878 338068 286906
rect 338132 286890 338160 287014
rect 337936 286816 337988 286822
rect 337936 286758 337988 286764
rect 337752 277374 337804 277380
rect 337842 277400 337898 277409
rect 337764 266665 337792 277374
rect 337842 277335 337898 277344
rect 337844 277296 337896 277302
rect 337844 277238 337896 277244
rect 337856 276865 337884 277238
rect 337842 276856 337898 276865
rect 337842 276791 337898 276800
rect 337844 276004 337896 276010
rect 337844 275946 337896 275952
rect 337856 275641 337884 275946
rect 337842 275632 337898 275641
rect 337842 275567 337898 275576
rect 337844 274644 337896 274650
rect 337844 274586 337896 274592
rect 337856 273737 337884 274586
rect 337842 273728 337898 273737
rect 337842 273663 337898 273672
rect 337844 273216 337896 273222
rect 337844 273158 337896 273164
rect 337856 272377 337884 273158
rect 337842 272368 337898 272377
rect 337842 272303 337898 272312
rect 337844 271856 337896 271862
rect 337844 271798 337896 271804
rect 337856 271153 337884 271798
rect 337842 271144 337898 271153
rect 337842 271079 337898 271088
rect 337844 270428 337896 270434
rect 337844 270370 337896 270376
rect 337856 269793 337884 270370
rect 337842 269784 337898 269793
rect 337842 269719 337898 269728
rect 337948 267345 337976 286758
rect 338040 278118 338068 286878
rect 338120 286884 338172 286890
rect 338120 286826 338172 286832
rect 338028 278112 338080 278118
rect 338028 278054 338080 278060
rect 338028 277976 338080 277982
rect 338028 277918 338080 277924
rect 338040 267889 338068 277918
rect 338026 267880 338082 267889
rect 338026 267815 338082 267824
rect 337934 267336 337990 267345
rect 337934 267271 337990 267280
rect 337750 266656 337806 266665
rect 337750 266591 337806 266600
rect 337658 265976 337714 265985
rect 337658 265911 337714 265920
rect 337566 264752 337622 264761
rect 337566 264687 337622 264696
rect 336830 264072 336886 264081
rect 336830 264007 336886 264016
rect 337474 263392 337530 263401
rect 337474 263327 337530 263336
rect 336832 262948 336884 262954
rect 336832 262890 336884 262896
rect 337384 262948 337436 262954
rect 337384 262890 337436 262896
rect 336096 256624 336148 256630
rect 336096 256566 336148 256572
rect 336004 84856 336056 84862
rect 336004 84798 336056 84804
rect 336108 3330 336136 256566
rect 336844 201414 336872 262890
rect 337016 262880 337068 262886
rect 337396 262857 337424 262890
rect 337488 262886 337516 263327
rect 337476 262880 337528 262886
rect 337016 262822 337068 262828
rect 337382 262848 337438 262857
rect 336924 259344 336976 259350
rect 336924 259286 336976 259292
rect 336936 258058 336964 259286
rect 336924 258052 336976 258058
rect 336924 257994 336976 258000
rect 336924 253224 336976 253230
rect 336924 253166 336976 253172
rect 336936 223582 336964 253166
rect 336924 223576 336976 223582
rect 336924 223518 336976 223524
rect 336832 201408 336884 201414
rect 336832 201350 336884 201356
rect 337028 201346 337056 262822
rect 337476 262822 337528 262828
rect 337382 262783 337438 262792
rect 337474 262168 337530 262177
rect 337474 262103 337530 262112
rect 337488 261526 337516 262103
rect 337660 261588 337712 261594
rect 337660 261530 337712 261536
rect 337476 261520 337528 261526
rect 337672 261497 337700 261530
rect 337476 261462 337528 261468
rect 337658 261488 337714 261497
rect 337658 261423 337714 261432
rect 337750 260808 337806 260817
rect 337750 260743 337806 260752
rect 337108 260296 337160 260302
rect 337108 260238 337160 260244
rect 337658 260264 337714 260273
rect 337120 259593 337148 260238
rect 337764 260234 337792 260743
rect 337658 260199 337714 260208
rect 337752 260228 337804 260234
rect 337672 260166 337700 260199
rect 337752 260170 337804 260176
rect 337660 260160 337712 260166
rect 337660 260102 337712 260108
rect 337106 259584 337162 259593
rect 337106 259519 337162 259528
rect 337120 253230 337148 259519
rect 337660 259412 337712 259418
rect 337660 259354 337712 259360
rect 337672 258369 337700 259354
rect 337658 258360 337714 258369
rect 337658 258295 337714 258304
rect 338776 258262 338804 289070
rect 339038 258632 339094 258641
rect 339038 258567 339094 258576
rect 338764 258256 338816 258262
rect 338764 258198 338816 258204
rect 339052 258058 339080 258567
rect 339040 258052 339092 258058
rect 339040 257994 339092 258000
rect 339420 255814 339448 575418
rect 360292 574048 360344 574054
rect 360292 573990 360344 573996
rect 426348 574048 426400 574054
rect 426348 573990 426400 573996
rect 351920 573980 351972 573986
rect 351920 573922 351972 573928
rect 349804 572688 349856 572694
rect 349804 572630 349856 572636
rect 341524 572620 341576 572626
rect 341524 572562 341576 572568
rect 340788 572144 340840 572150
rect 340788 572086 340840 572092
rect 340800 397882 340828 572086
rect 340880 453416 340932 453422
rect 340880 453358 340932 453364
rect 340892 422294 340920 453358
rect 340892 422266 341104 422294
rect 340492 397854 340828 397882
rect 341076 397882 341104 422266
rect 341536 401538 341564 572562
rect 345020 572552 345072 572558
rect 345020 572494 345072 572500
rect 342904 453348 342956 453354
rect 342904 453290 342956 453296
rect 342260 409352 342312 409358
rect 342260 409294 342312 409300
rect 341524 401532 341576 401538
rect 341524 401474 341576 401480
rect 342272 397882 342300 409294
rect 342916 401266 342944 453290
rect 345032 422294 345060 572494
rect 345032 422266 345336 422294
rect 342904 401260 342956 401266
rect 342904 401202 342956 401208
rect 343916 401056 343968 401062
rect 343916 400998 343968 401004
rect 343928 397882 343956 400998
rect 344744 400852 344796 400858
rect 344744 400794 344796 400800
rect 344756 397882 344784 400794
rect 341076 397854 341504 397882
rect 342272 397854 342516 397882
rect 343620 397854 343956 397882
rect 344632 397854 344784 397882
rect 345308 397882 345336 422266
rect 349436 406020 349488 406026
rect 349436 405962 349488 405968
rect 349068 401600 349120 401606
rect 349068 401542 349120 401548
rect 347872 401532 347924 401538
rect 347872 401474 347924 401480
rect 346400 401260 346452 401266
rect 346400 401202 346452 401208
rect 346412 397882 346440 401202
rect 345308 397854 345736 397882
rect 346412 397854 346748 397882
rect 347884 397746 347912 401474
rect 349080 397882 349108 401542
rect 348864 397854 349108 397882
rect 349448 397882 349476 405962
rect 349816 400790 349844 572630
rect 350632 401124 350684 401130
rect 350632 401066 350684 401072
rect 349804 400784 349856 400790
rect 349804 400726 349856 400732
rect 350644 397882 350672 401066
rect 351932 398154 351960 573922
rect 357440 573300 357492 573306
rect 357440 573242 357492 573248
rect 356060 572484 356112 572490
rect 356060 572426 356112 572432
rect 353944 456204 353996 456210
rect 353944 456146 353996 456152
rect 353668 406088 353720 406094
rect 353668 406030 353720 406036
rect 353208 401532 353260 401538
rect 353208 401474 353260 401480
rect 351932 398126 352006 398154
rect 349448 397854 349876 397882
rect 350644 397854 350980 397882
rect 351978 397868 352006 398126
rect 353220 397882 353248 401474
rect 353096 397854 353248 397882
rect 353680 397882 353708 406030
rect 353956 401266 353984 456146
rect 356072 422294 356100 572426
rect 357452 422294 357480 573242
rect 360304 422294 360332 573990
rect 367008 573980 367060 573986
rect 367008 573922 367060 573928
rect 363604 573232 363656 573238
rect 363604 573174 363656 573180
rect 356072 422266 356928 422294
rect 357452 422266 357940 422294
rect 360304 422266 361068 422294
rect 353944 401260 353996 401266
rect 353944 401202 353996 401208
rect 354956 401192 355008 401198
rect 354956 401134 355008 401140
rect 354968 397882 354996 401134
rect 356520 401124 356572 401130
rect 356520 401066 356572 401072
rect 356532 397882 356560 401066
rect 353680 397854 354108 397882
rect 354968 397854 355212 397882
rect 356224 397854 356560 397882
rect 356900 397882 356928 422266
rect 357912 397882 357940 422266
rect 360200 401260 360252 401266
rect 360200 401202 360252 401208
rect 359648 400648 359700 400654
rect 359648 400590 359700 400596
rect 359660 397882 359688 400590
rect 356900 397854 357328 397882
rect 357912 397854 358340 397882
rect 359352 397854 359688 397882
rect 360212 397882 360240 401202
rect 361040 397882 361068 422266
rect 362868 401260 362920 401266
rect 362868 401202 362920 401208
rect 362880 397882 362908 401202
rect 363616 400790 363644 573174
rect 364984 410508 365036 410514
rect 364984 410450 365036 410456
rect 363236 400784 363288 400790
rect 363236 400726 363288 400732
rect 363604 400784 363656 400790
rect 363604 400726 363656 400732
rect 360212 397854 360456 397882
rect 361040 397854 361468 397882
rect 362572 397854 362908 397882
rect 363248 397882 363276 400726
rect 364524 400716 364576 400722
rect 364524 400658 364576 400664
rect 364536 397882 364564 400658
rect 364996 400314 365024 410450
rect 364984 400308 365036 400314
rect 364984 400250 365036 400256
rect 366456 400308 366508 400314
rect 366456 400250 366508 400256
rect 365996 400240 366048 400246
rect 365996 400182 366048 400188
rect 366008 397882 366036 400182
rect 363248 397854 363584 397882
rect 364536 397854 364688 397882
rect 365700 397854 366036 397882
rect 366468 397882 366496 400250
rect 367020 400246 367048 573922
rect 367100 573912 367152 573918
rect 367100 573854 367152 573860
rect 369768 573912 369820 573918
rect 369768 573854 369820 573860
rect 367112 422294 367140 573854
rect 367112 422266 367416 422294
rect 367008 400240 367060 400246
rect 367008 400182 367060 400188
rect 367388 397882 367416 422266
rect 369780 400246 369808 573854
rect 395344 573844 395396 573850
rect 395344 573786 395396 573792
rect 407028 573844 407080 573850
rect 407028 573786 407080 573792
rect 370504 572416 370556 572422
rect 370504 572358 370556 572364
rect 382188 572416 382240 572422
rect 382188 572358 382240 572364
rect 369952 411256 370004 411262
rect 369952 411198 370004 411204
rect 369124 400240 369176 400246
rect 369124 400182 369176 400188
rect 369768 400240 369820 400246
rect 369768 400182 369820 400188
rect 369136 397882 369164 400182
rect 369964 397882 369992 411198
rect 370516 400654 370544 572358
rect 374644 572348 374696 572354
rect 374644 572290 374696 572296
rect 379428 572348 379480 572354
rect 379428 572290 379480 572296
rect 371884 411188 371936 411194
rect 371884 411130 371936 411136
rect 370596 401464 370648 401470
rect 370596 401406 370648 401412
rect 370504 400648 370556 400654
rect 370504 400590 370556 400596
rect 366468 397854 366804 397882
rect 367388 397854 367816 397882
rect 368828 397854 369164 397882
rect 369932 397854 369992 397882
rect 370608 397882 370636 401406
rect 371896 400246 371924 411130
rect 374000 409216 374052 409222
rect 374000 409158 374052 409164
rect 372344 400716 372396 400722
rect 372344 400658 372396 400664
rect 371884 400240 371936 400246
rect 371884 400182 371936 400188
rect 372356 397882 372384 400658
rect 372712 400240 372764 400246
rect 372712 400182 372764 400188
rect 370608 397854 370944 397882
rect 372048 397854 372384 397882
rect 372724 397882 372752 400182
rect 374012 397882 374040 409158
rect 374656 400246 374684 572290
rect 378968 411120 379020 411126
rect 378968 411062 379020 411068
rect 376852 409284 376904 409290
rect 376852 409226 376904 409232
rect 375288 402280 375340 402286
rect 375288 402222 375340 402228
rect 374644 400240 374696 400246
rect 374644 400182 374696 400188
rect 375300 397882 375328 402222
rect 375932 400240 375984 400246
rect 375932 400182 375984 400188
rect 372724 397854 373060 397882
rect 374012 397854 374164 397882
rect 375176 397854 375328 397882
rect 375944 397882 375972 400182
rect 376864 397882 376892 409226
rect 378600 400240 378652 400246
rect 378600 400182 378652 400188
rect 378612 397882 378640 400182
rect 375944 397854 376280 397882
rect 376864 397854 377292 397882
rect 378304 397854 378640 397882
rect 378980 397882 379008 411062
rect 379440 400246 379468 572290
rect 379980 409148 380032 409154
rect 379980 409090 380032 409096
rect 379428 400240 379480 400246
rect 379428 400182 379480 400188
rect 379992 397882 380020 409090
rect 382200 402974 382228 572358
rect 388444 572280 388496 572286
rect 388444 572222 388496 572228
rect 382924 572076 382976 572082
rect 382924 572018 382976 572024
rect 381924 402946 382228 402974
rect 381924 397882 381952 402946
rect 382936 400722 382964 572018
rect 387800 456136 387852 456142
rect 387800 456078 387852 456084
rect 387812 422294 387840 456078
rect 387812 422266 388392 422294
rect 385316 411052 385368 411058
rect 385316 410994 385368 411000
rect 383660 410644 383712 410650
rect 383660 410586 383712 410592
rect 382924 400716 382976 400722
rect 382924 400658 382976 400664
rect 382280 400648 382332 400654
rect 382280 400590 382332 400596
rect 378980 397854 379408 397882
rect 379992 397854 380420 397882
rect 381524 397854 381952 397882
rect 382292 397882 382320 400590
rect 383672 397882 383700 410586
rect 384948 402348 385000 402354
rect 384948 402290 385000 402296
rect 384960 397882 384988 402290
rect 382292 397854 382536 397882
rect 383640 397854 383700 397882
rect 384652 397854 384988 397882
rect 385328 397882 385356 410994
rect 386420 410576 386472 410582
rect 386420 410518 386472 410524
rect 386432 397882 386460 410518
rect 388076 402416 388128 402422
rect 388076 402358 388128 402364
rect 388088 397882 388116 402358
rect 385328 397854 385756 397882
rect 386432 397854 386768 397882
rect 387780 397854 388116 397882
rect 388364 397882 388392 422266
rect 388456 400246 388484 572222
rect 393964 572008 394016 572014
rect 393964 571950 394016 571956
rect 389456 412208 389508 412214
rect 389456 412150 389508 412156
rect 388444 400240 388496 400246
rect 388444 400182 388496 400188
rect 389468 397882 389496 412150
rect 392676 412140 392728 412146
rect 392676 412082 392728 412088
rect 391296 402484 391348 402490
rect 391296 402426 391348 402432
rect 391308 397882 391336 402426
rect 392032 400240 392084 400246
rect 392032 400182 392084 400188
rect 388364 397854 388884 397882
rect 389468 397854 389896 397882
rect 391000 397854 391336 397882
rect 392044 397746 392072 400182
rect 392688 397882 392716 412082
rect 393976 400314 394004 571950
rect 394792 410984 394844 410990
rect 394792 410926 394844 410932
rect 394424 403640 394476 403646
rect 394424 403582 394476 403588
rect 393964 400308 394016 400314
rect 393964 400250 394016 400256
rect 394436 397882 394464 403582
rect 392688 397854 393116 397882
rect 394128 397854 394464 397882
rect 394804 397882 394832 410926
rect 395356 400654 395384 573786
rect 399484 573776 399536 573782
rect 399484 573718 399536 573724
rect 404268 573776 404320 573782
rect 404268 573718 404320 573724
rect 396724 572212 396776 572218
rect 396724 572154 396776 572160
rect 396080 412072 396132 412078
rect 396080 412014 396132 412020
rect 395344 400648 395396 400654
rect 395344 400590 395396 400596
rect 396092 397882 396120 412014
rect 396736 400246 396764 572154
rect 398932 412004 398984 412010
rect 398932 411946 398984 411952
rect 397368 403708 397420 403714
rect 397368 403650 397420 403656
rect 396724 400240 396776 400246
rect 396724 400182 396776 400188
rect 397380 397882 397408 403650
rect 398012 400240 398064 400246
rect 398012 400182 398064 400188
rect 394804 397854 395232 397882
rect 396092 397854 396244 397882
rect 397256 397854 397408 397882
rect 398024 397882 398052 400182
rect 398944 397882 398972 411946
rect 399496 400518 399524 573718
rect 400220 456068 400272 456074
rect 400220 456010 400272 456016
rect 400232 422294 400260 456010
rect 400232 422266 401088 422294
rect 400772 402552 400824 402558
rect 400772 402494 400824 402500
rect 399484 400512 399536 400518
rect 399484 400454 399536 400460
rect 400784 397882 400812 402494
rect 398024 397854 398360 397882
rect 398944 397854 399372 397882
rect 400476 397854 400812 397882
rect 401060 397882 401088 422266
rect 403624 410916 403676 410922
rect 403624 410858 403676 410864
rect 402244 400308 402296 400314
rect 402244 400250 402296 400256
rect 402256 397882 402284 400250
rect 403636 400246 403664 410858
rect 404280 402974 404308 573718
rect 405740 411936 405792 411942
rect 405740 411878 405792 411884
rect 404004 402946 404308 402974
rect 403624 400240 403676 400246
rect 403624 400182 403676 400188
rect 404004 397882 404032 402946
rect 404360 400240 404412 400246
rect 404360 400182 404412 400188
rect 401060 397854 401488 397882
rect 402256 397854 402592 397882
rect 403604 397854 404032 397882
rect 404372 397882 404400 400182
rect 405752 397882 405780 411878
rect 407040 397882 407068 573786
rect 410524 573708 410576 573714
rect 410524 573650 410576 573656
rect 416688 573708 416740 573714
rect 416688 573650 416740 573656
rect 407764 573640 407816 573646
rect 407764 573582 407816 573588
rect 407396 410780 407448 410786
rect 407396 410722 407448 410728
rect 404372 397854 404708 397882
rect 405720 397854 405780 397882
rect 406732 397854 407068 397882
rect 407408 397882 407436 410722
rect 407776 400382 407804 573582
rect 409144 573028 409196 573034
rect 409144 572970 409196 572976
rect 409156 400858 409184 572970
rect 410536 422294 410564 573650
rect 411904 573640 411956 573646
rect 411904 573582 411956 573588
rect 410536 422266 410656 422294
rect 410432 410848 410484 410854
rect 410432 410790 410484 410796
rect 410444 402974 410472 410790
rect 410444 402946 410564 402974
rect 409144 400852 409196 400858
rect 409144 400794 409196 400800
rect 408500 400716 408552 400722
rect 408500 400658 408552 400664
rect 407764 400376 407816 400382
rect 407764 400318 407816 400324
rect 408512 397882 408540 400658
rect 410248 400240 410300 400246
rect 410248 400182 410300 400188
rect 410260 397882 410288 400182
rect 407408 397854 407836 397882
rect 408512 397854 408848 397882
rect 409952 397854 410288 397882
rect 410536 397882 410564 402946
rect 410628 400858 410656 422266
rect 410616 400852 410668 400858
rect 410616 400794 410668 400800
rect 411720 400512 411772 400518
rect 411720 400454 411772 400460
rect 411732 397882 411760 400454
rect 411916 400246 411944 573582
rect 413284 573504 413336 573510
rect 413284 573446 413336 573452
rect 414664 573504 414716 573510
rect 414664 573446 414716 573452
rect 413296 400518 413324 573446
rect 414112 410712 414164 410718
rect 414112 410654 414164 410660
rect 413284 400512 413336 400518
rect 413284 400454 413336 400460
rect 411904 400240 411956 400246
rect 411904 400182 411956 400188
rect 413376 400240 413428 400246
rect 413376 400182 413428 400188
rect 413388 397882 413416 400182
rect 414124 398154 414152 410654
rect 414676 400246 414704 573446
rect 416700 402974 416728 573650
rect 417424 573572 417476 573578
rect 417424 573514 417476 573520
rect 419448 573572 419500 573578
rect 419448 573514 419500 573520
rect 416872 406156 416924 406162
rect 416872 406098 416924 406104
rect 416608 402946 416728 402974
rect 414848 400648 414900 400654
rect 414848 400590 414900 400596
rect 414664 400240 414716 400246
rect 414664 400182 414716 400188
rect 414124 398126 414198 398154
rect 410536 397854 410964 397882
rect 411732 397854 412068 397882
rect 413080 397854 413416 397882
rect 414170 397868 414198 398126
rect 414860 397882 414888 400590
rect 416608 397882 416636 402946
rect 414860 397854 415196 397882
rect 416208 397854 416636 397882
rect 416884 397882 416912 406098
rect 417436 400722 417464 573514
rect 418160 400784 418212 400790
rect 418160 400726 418212 400732
rect 417424 400716 417476 400722
rect 417424 400658 417476 400664
rect 418172 397882 418200 400726
rect 419460 397882 419488 573514
rect 421564 573436 421616 573442
rect 421564 573378 421616 573384
rect 423588 573436 423640 573442
rect 423588 573378 423640 573384
rect 420184 572960 420236 572966
rect 420184 572902 420236 572908
rect 420000 406224 420052 406230
rect 420000 406166 420052 406172
rect 416884 397854 417312 397882
rect 418172 397854 418324 397882
rect 419428 397854 419488 397882
rect 420012 397882 420040 406166
rect 420196 401606 420224 572902
rect 421576 401606 421604 573378
rect 420184 401600 420236 401606
rect 420184 401542 420236 401548
rect 421564 401600 421616 401606
rect 421564 401542 421616 401548
rect 421196 400376 421248 400382
rect 421196 400318 421248 400324
rect 421208 397882 421236 400318
rect 423600 400246 423628 573378
rect 423772 406292 423824 406298
rect 423772 406234 423824 406240
rect 422852 400240 422904 400246
rect 422852 400182 422904 400188
rect 423588 400240 423640 400246
rect 423588 400182 423640 400188
rect 422864 397882 422892 400182
rect 423784 397882 423812 406234
rect 426360 402974 426388 573990
rect 431224 573368 431276 573374
rect 431224 573310 431276 573316
rect 433248 573368 433300 573374
rect 433248 573310 433300 573316
rect 429108 573300 429160 573306
rect 429108 573242 429160 573248
rect 426440 406360 426492 406366
rect 426440 406302 426492 406308
rect 426084 402946 426388 402974
rect 424324 400512 424376 400518
rect 424324 400454 424376 400460
rect 420012 397854 420440 397882
rect 421208 397854 421544 397882
rect 422556 397854 422892 397882
rect 423660 397854 423812 397882
rect 424336 397882 424364 400454
rect 426084 397882 426112 402946
rect 424336 397854 424672 397882
rect 425684 397854 426112 397882
rect 426452 397882 426480 406302
rect 427820 400852 427872 400858
rect 427820 400794 427872 400800
rect 427832 397882 427860 400794
rect 429120 397882 429148 573242
rect 429476 407108 429528 407114
rect 429476 407050 429528 407056
rect 426452 397854 426788 397882
rect 427800 397854 427860 397882
rect 428904 397854 429148 397882
rect 429488 397882 429516 407050
rect 431236 400858 431264 573310
rect 432696 407040 432748 407046
rect 432696 406982 432748 406988
rect 431224 400852 431276 400858
rect 431224 400794 431276 400800
rect 430672 400716 430724 400722
rect 430672 400658 430724 400664
rect 430684 397882 430712 400658
rect 432328 400240 432380 400246
rect 432328 400182 432380 400188
rect 432340 397882 432368 400182
rect 429488 397854 429916 397882
rect 430684 397854 431020 397882
rect 432032 397854 432368 397882
rect 432708 397882 432736 406982
rect 433260 400246 433288 573310
rect 436008 573232 436060 573238
rect 436008 573174 436060 573180
rect 433800 401600 433852 401606
rect 433800 401542 433852 401548
rect 433248 400240 433300 400246
rect 433248 400182 433300 400188
rect 433812 397882 433840 401542
rect 436020 400246 436048 573174
rect 438768 573164 438820 573170
rect 438768 573106 438820 573112
rect 436192 406972 436244 406978
rect 436192 406914 436244 406920
rect 435456 400240 435508 400246
rect 435456 400182 435508 400188
rect 436008 400240 436060 400246
rect 436008 400182 436060 400188
rect 435468 397882 435496 400182
rect 436204 398154 436232 406914
rect 436928 400852 436980 400858
rect 436928 400794 436980 400800
rect 436204 398126 436278 398154
rect 432708 397854 433136 397882
rect 433812 397854 434148 397882
rect 435160 397854 435496 397882
rect 436250 397868 436278 398126
rect 436940 397882 436968 400794
rect 438780 397882 438808 573106
rect 441528 573096 441580 573102
rect 441528 573038 441580 573044
rect 438952 406904 439004 406910
rect 438952 406846 439004 406852
rect 436940 397854 437276 397882
rect 438380 397854 438808 397882
rect 438964 397882 438992 406846
rect 440240 401396 440292 401402
rect 440240 401338 440292 401344
rect 440252 397882 440280 401338
rect 441540 397882 441568 573038
rect 443644 572892 443696 572898
rect 443644 572834 443696 572840
rect 442172 406836 442224 406842
rect 442172 406778 442224 406784
rect 438964 397854 439392 397882
rect 440252 397854 440496 397882
rect 441508 397854 441568 397882
rect 442184 397882 442212 406778
rect 443656 401606 443684 572834
rect 443644 401600 443696 401606
rect 443644 401542 443696 401548
rect 443276 401328 443328 401334
rect 443276 401270 443328 401276
rect 443288 397882 443316 401270
rect 444392 397882 444420 577594
rect 447152 422294 447180 601666
rect 447152 422266 447456 422294
rect 447048 401396 447100 401402
rect 447048 401338 447100 401344
rect 446036 401328 446088 401334
rect 446036 401270 446088 401276
rect 446048 397882 446076 401270
rect 447060 397882 447088 401338
rect 442184 397854 442612 397882
rect 443288 397854 443624 397882
rect 444392 397854 444636 397882
rect 445740 397854 446076 397882
rect 446752 397854 447088 397882
rect 447428 397882 447456 422266
rect 449164 401532 449216 401538
rect 449164 401474 449216 401480
rect 449176 397882 449204 401474
rect 449912 398154 449940 609962
rect 451292 422294 451320 618870
rect 452212 618322 452240 618870
rect 452200 618316 452252 618322
rect 452200 618258 452252 618264
rect 451292 422266 451688 422294
rect 451096 401600 451148 401606
rect 451096 401542 451148 401548
rect 449912 398126 449986 398154
rect 447428 397854 447856 397882
rect 448868 397854 449204 397882
rect 449958 397868 449986 398126
rect 451108 397882 451136 401542
rect 450984 397854 451136 397882
rect 451660 397882 451688 422266
rect 453396 400852 453448 400858
rect 453396 400794 453448 400800
rect 453408 397882 453436 400794
rect 454052 398154 454080 626554
rect 454052 398126 454126 398154
rect 451660 397854 452088 397882
rect 453100 397854 453436 397882
rect 454098 397868 454126 398126
rect 455340 397882 455368 680342
rect 459468 585200 459520 585206
rect 459468 585142 459520 585148
rect 459008 409420 459060 409426
rect 459008 409362 459060 409368
rect 455880 400988 455932 400994
rect 455880 400930 455932 400936
rect 455216 397854 455368 397882
rect 455892 397882 455920 400930
rect 456984 400920 457036 400926
rect 456984 400862 457036 400868
rect 456996 397882 457024 400862
rect 458640 400240 458692 400246
rect 458640 400182 458692 400188
rect 458652 397882 458680 400182
rect 455892 397854 456228 397882
rect 456996 397854 457332 397882
rect 458344 397854 458680 397882
rect 459020 397882 459048 409362
rect 459480 400246 459508 585142
rect 460952 422294 460980 700334
rect 462240 700210 462268 700470
rect 462332 700330 462360 703520
rect 472072 701004 472124 701010
rect 472072 700946 472124 700952
rect 469220 700936 469272 700942
rect 469220 700878 469272 700884
rect 467932 700800 467984 700806
rect 467932 700742 467984 700748
rect 467840 700732 467892 700738
rect 467840 700674 467892 700680
rect 465080 700664 465132 700670
rect 465080 700606 465132 700612
rect 463700 700460 463752 700466
rect 463700 700402 463752 700408
rect 462412 700392 462464 700398
rect 462412 700334 462464 700340
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 462240 700182 462360 700210
rect 460952 422266 461164 422294
rect 460018 409184 460074 409193
rect 460018 409119 460074 409128
rect 459468 400240 459520 400246
rect 459468 400182 459520 400188
rect 460032 397882 460060 409119
rect 461136 397882 461164 422266
rect 462332 400178 462360 700182
rect 462320 400172 462372 400178
rect 462320 400114 462372 400120
rect 462424 397882 462452 700334
rect 463712 422294 463740 700402
rect 465092 422294 465120 700606
rect 466460 700596 466512 700602
rect 466460 700538 466512 700544
rect 463712 422266 464292 422294
rect 465092 422266 465304 422294
rect 463240 400172 463292 400178
rect 463240 400114 463292 400120
rect 463252 397882 463280 400114
rect 464264 397882 464292 422266
rect 465276 397882 465304 422266
rect 466472 397882 466500 700538
rect 467852 400178 467880 700674
rect 467840 400172 467892 400178
rect 467840 400114 467892 400120
rect 467944 397882 467972 700742
rect 469232 422294 469260 700878
rect 470600 700868 470652 700874
rect 470600 700810 470652 700816
rect 469232 422266 469536 422294
rect 468576 400172 468628 400178
rect 468576 400114 468628 400120
rect 459020 397854 459448 397882
rect 460032 397854 460460 397882
rect 461136 397854 461564 397882
rect 462424 397854 462576 397882
rect 463252 397854 463588 397882
rect 464264 397854 464692 397882
rect 465276 397854 465704 397882
rect 466472 397854 466808 397882
rect 467820 397854 467972 397882
rect 468588 397882 468616 400114
rect 469508 397882 469536 422266
rect 470612 397882 470640 700810
rect 471980 700256 472032 700262
rect 471980 700198 472032 700204
rect 471992 398018 472020 700198
rect 472084 398154 472112 700946
rect 472808 700324 472860 700330
rect 472808 700266 472860 700272
rect 472716 700188 472768 700194
rect 472716 700130 472768 700136
rect 472622 627736 472678 627745
rect 472622 627671 472678 627680
rect 472636 626618 472664 627671
rect 472624 626612 472676 626618
rect 472624 626554 472676 626560
rect 472530 623520 472586 623529
rect 472530 623455 472586 623464
rect 472544 623082 472572 623455
rect 472164 623076 472216 623082
rect 472164 623018 472216 623024
rect 472532 623076 472584 623082
rect 472532 623018 472584 623024
rect 472176 400858 472204 623018
rect 472622 619440 472678 619449
rect 472622 619375 472678 619384
rect 472636 618322 472664 619375
rect 472624 618316 472676 618322
rect 472624 618258 472676 618264
rect 472530 615224 472586 615233
rect 472530 615159 472586 615168
rect 472544 614786 472572 615159
rect 472256 614780 472308 614786
rect 472256 614722 472308 614728
rect 472532 614780 472584 614786
rect 472532 614722 472584 614728
rect 472268 401606 472296 614722
rect 472622 611144 472678 611153
rect 472622 611079 472678 611088
rect 472636 610026 472664 611079
rect 472624 610020 472676 610026
rect 472624 609962 472676 609968
rect 472438 606928 472494 606937
rect 472438 606863 472494 606872
rect 472452 606490 472480 606863
rect 472440 606484 472492 606490
rect 472440 606426 472492 606432
rect 472452 586514 472480 606426
rect 472622 602848 472678 602857
rect 472622 602783 472678 602792
rect 472636 601730 472664 602783
rect 472624 601724 472676 601730
rect 472624 601666 472676 601672
rect 472622 590336 472678 590345
rect 472622 590271 472678 590280
rect 472636 589354 472664 590271
rect 472624 589348 472676 589354
rect 472624 589290 472676 589296
rect 472360 586486 472480 586514
rect 472256 401600 472308 401606
rect 472256 401542 472308 401548
rect 472360 401402 472388 586486
rect 472622 586256 472678 586265
rect 472622 586191 472678 586200
rect 472636 585206 472664 586191
rect 472624 585200 472676 585206
rect 472624 585142 472676 585148
rect 472532 578196 472584 578202
rect 472532 578138 472584 578144
rect 472440 578128 472492 578134
rect 472440 578070 472492 578076
rect 472452 577590 472480 578070
rect 472544 577862 472572 578138
rect 472622 577960 472678 577969
rect 472622 577895 472678 577904
rect 472532 577856 472584 577862
rect 472532 577798 472584 577804
rect 472440 577584 472492 577590
rect 472440 577526 472492 577532
rect 472348 401396 472400 401402
rect 472348 401338 472400 401344
rect 472452 400994 472480 577526
rect 472544 401334 472572 577798
rect 472636 577522 472664 577895
rect 472624 577516 472676 577522
rect 472624 577458 472676 577464
rect 472532 401328 472584 401334
rect 472532 401270 472584 401276
rect 472440 400988 472492 400994
rect 472440 400930 472492 400936
rect 472164 400852 472216 400858
rect 472164 400794 472216 400800
rect 472728 400314 472756 700130
rect 472820 400382 472848 700266
rect 472900 700120 472952 700126
rect 472900 700062 472952 700068
rect 472808 400376 472860 400382
rect 472808 400318 472860 400324
rect 472716 400308 472768 400314
rect 472716 400250 472768 400256
rect 472912 400246 472940 700062
rect 478524 699718 478552 703520
rect 491300 700052 491352 700058
rect 491300 699994 491352 700000
rect 475384 699712 475436 699718
rect 475384 699654 475436 699660
rect 478512 699712 478564 699718
rect 478512 699654 478564 699660
rect 472990 598632 473046 598641
rect 472990 598567 473046 598576
rect 473004 578202 473032 598567
rect 473082 594552 473138 594561
rect 473082 594487 473138 594496
rect 472992 578196 473044 578202
rect 472992 578138 473044 578144
rect 473096 578134 473124 594487
rect 473174 582040 473230 582049
rect 473174 581975 473230 581984
rect 473084 578128 473136 578134
rect 473084 578070 473136 578076
rect 473188 575482 473216 581975
rect 475396 576162 475424 699654
rect 491312 692774 491340 699994
rect 491312 692746 491708 692774
rect 483478 680640 483534 680649
rect 483478 680575 483534 680584
rect 483492 680406 483520 680575
rect 483480 680400 483532 680406
rect 483480 680342 483532 680348
rect 491680 680082 491708 692746
rect 511000 683114 511028 703520
rect 527192 699718 527220 703520
rect 543476 700330 543504 703520
rect 530584 700324 530636 700330
rect 530584 700266 530636 700272
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 528560 699712 528612 699718
rect 528560 699654 528612 699660
rect 510908 683086 511028 683114
rect 491680 680054 492108 680082
rect 487264 676314 487600 676342
rect 490668 676314 491004 676342
rect 482928 674212 482980 674218
rect 482928 674154 482980 674160
rect 477408 674144 477460 674150
rect 477408 674086 477460 674092
rect 477420 629762 477448 674086
rect 482940 632126 482968 674154
rect 487264 674150 487292 676314
rect 490668 674218 490696 676314
rect 490656 674212 490708 674218
rect 490656 674154 490708 674160
rect 487252 674144 487304 674150
rect 487252 674086 487304 674092
rect 491680 663794 491708 680054
rect 494440 676314 494776 676342
rect 494440 673946 494468 676314
rect 493324 673940 493376 673946
rect 493324 673882 493376 673888
rect 494428 673940 494480 673946
rect 494428 673882 494480 673888
rect 491588 663766 491708 663794
rect 491588 632398 491616 663766
rect 486884 632392 486936 632398
rect 486884 632334 486936 632340
rect 491576 632392 491628 632398
rect 491576 632334 491628 632340
rect 482008 632120 482060 632126
rect 482008 632062 482060 632068
rect 482928 632120 482980 632126
rect 482928 632062 482980 632068
rect 477158 629734 477448 629762
rect 482020 629748 482048 632062
rect 486896 629748 486924 632334
rect 493336 632126 493364 673882
rect 491852 632120 491904 632126
rect 491852 632062 491904 632068
rect 493324 632120 493376 632126
rect 496832 632074 496860 680068
rect 499592 680054 500342 680082
rect 502444 680054 502872 680082
rect 506492 680054 507380 680082
rect 499500 673538 499528 676328
rect 499488 673532 499540 673538
rect 499488 673474 499540 673480
rect 499592 632194 499620 680054
rect 501998 676314 502288 676342
rect 500224 673532 500276 673538
rect 500224 673474 500276 673480
rect 499580 632188 499632 632194
rect 499580 632130 499632 632136
rect 500236 632126 500264 673474
rect 502260 632942 502288 676314
rect 502248 632936 502300 632942
rect 502248 632878 502300 632884
rect 502444 632874 502472 680054
rect 505572 674354 505600 676328
rect 505560 674348 505612 674354
rect 505560 674290 505612 674296
rect 506388 674348 506440 674354
rect 506388 674290 506440 674296
rect 502432 632868 502484 632874
rect 502432 632810 502484 632816
rect 506400 632806 506428 674290
rect 506388 632800 506440 632806
rect 506388 632742 506440 632748
rect 506492 632738 506520 680054
rect 510908 679221 510936 683086
rect 510894 679212 510950 679221
rect 510894 679147 510950 679156
rect 511448 632936 511500 632942
rect 511448 632878 511500 632884
rect 506480 632732 506532 632738
rect 506480 632674 506532 632680
rect 506572 632188 506624 632194
rect 506572 632130 506624 632136
rect 493324 632062 493376 632068
rect 491864 629748 491892 632062
rect 496740 632046 496860 632074
rect 500224 632120 500276 632126
rect 500224 632062 500276 632068
rect 501604 632120 501656 632126
rect 501604 632062 501656 632068
rect 496740 629748 496768 632046
rect 501616 629748 501644 632062
rect 506584 629748 506612 632130
rect 511460 629748 511488 632878
rect 516324 632868 516376 632874
rect 516324 632810 516376 632816
rect 516336 629748 516364 632810
rect 521292 632800 521344 632806
rect 521292 632742 521344 632748
rect 521304 629748 521332 632742
rect 526168 632732 526220 632738
rect 526168 632674 526220 632680
rect 526180 629748 526208 632674
rect 528572 576162 528600 699654
rect 529204 683188 529256 683194
rect 529204 683130 529256 683136
rect 475384 576156 475436 576162
rect 475384 576098 475436 576104
rect 480168 576156 480220 576162
rect 480168 576098 480220 576104
rect 528560 576156 528612 576162
rect 528560 576098 528612 576104
rect 474752 576014 475502 576042
rect 473176 575476 473228 575482
rect 473176 575418 473228 575424
rect 474752 401062 474780 576014
rect 475384 575884 475436 575890
rect 475384 575826 475436 575832
rect 474740 401056 474792 401062
rect 474740 400998 474792 401004
rect 474832 400308 474884 400314
rect 474832 400250 474884 400256
rect 472900 400240 472952 400246
rect 472900 400182 472952 400188
rect 473820 400240 473872 400246
rect 473820 400182 473872 400188
rect 472084 398126 472664 398154
rect 471992 397990 472066 398018
rect 468588 397854 468924 397882
rect 469508 397854 469936 397882
rect 470612 397854 471040 397882
rect 472038 397868 472066 397990
rect 472636 397882 472664 398126
rect 473832 397882 473860 400182
rect 474844 397882 474872 400250
rect 475396 400246 475424 575826
rect 476764 572824 476816 572830
rect 476764 572766 476816 572772
rect 476776 401130 476804 572766
rect 477052 572150 477080 575892
rect 478708 573034 478736 575892
rect 478696 573028 478748 573034
rect 478696 572970 478748 572976
rect 478144 572756 478196 572762
rect 478144 572698 478196 572704
rect 477040 572144 477092 572150
rect 477040 572086 477092 572092
rect 478156 401198 478184 572698
rect 478144 401192 478196 401198
rect 478144 401134 478196 401140
rect 476764 401124 476816 401130
rect 476764 401066 476816 401072
rect 478696 400920 478748 400926
rect 478696 400862 478748 400868
rect 476948 400376 477000 400382
rect 476948 400318 477000 400324
rect 475384 400240 475436 400246
rect 475384 400182 475436 400188
rect 476120 400240 476172 400246
rect 476120 400182 476172 400188
rect 476132 397882 476160 400182
rect 476960 397882 476988 400318
rect 478708 397882 478736 400862
rect 480180 400246 480208 576098
rect 480364 572966 480392 575892
rect 480352 572960 480404 572966
rect 480352 572902 480404 572908
rect 482020 572898 482048 575892
rect 482284 573028 482336 573034
rect 482284 572970 482336 572976
rect 482008 572892 482060 572898
rect 482008 572834 482060 572840
rect 480904 572756 480956 572762
rect 480904 572698 480956 572704
rect 480916 401266 480944 572698
rect 482296 401470 482324 572970
rect 483584 572830 483612 575892
rect 485240 572966 485268 575892
rect 485228 572960 485280 572966
rect 485228 572902 485280 572908
rect 483572 572824 483624 572830
rect 483572 572766 483624 572772
rect 486896 572762 486924 575892
rect 488552 573986 488580 575892
rect 488540 573980 488592 573986
rect 488540 573922 488592 573928
rect 490208 573918 490236 575892
rect 490196 573912 490248 573918
rect 490196 573854 490248 573860
rect 491772 573034 491800 575892
rect 492692 575878 493442 575906
rect 491760 573028 491812 573034
rect 491760 572970 491812 572976
rect 486884 572756 486936 572762
rect 486884 572698 486936 572704
rect 482376 536852 482428 536858
rect 482376 536794 482428 536800
rect 482284 401464 482336 401470
rect 482284 401406 482336 401412
rect 480904 401260 480956 401266
rect 480904 401202 480956 401208
rect 479708 400240 479760 400246
rect 479708 400182 479760 400188
rect 480168 400240 480220 400246
rect 480168 400182 480220 400188
rect 479720 397882 479748 400182
rect 472636 397854 473064 397882
rect 473832 397854 474168 397882
rect 474844 397854 475180 397882
rect 476132 397854 476284 397882
rect 476960 397854 477296 397882
rect 478400 397854 478736 397882
rect 479412 397854 479748 397882
rect 347852 397718 347912 397746
rect 392012 397718 392072 397746
rect 482008 382220 482060 382226
rect 482008 382162 482060 382168
rect 482020 381585 482048 382162
rect 482006 381576 482062 381585
rect 482006 381511 482062 381520
rect 482192 378208 482244 378214
rect 482192 378150 482244 378156
rect 482204 373994 482232 378150
rect 482284 378140 482336 378146
rect 482284 378082 482336 378088
rect 482296 376961 482324 378082
rect 482282 376952 482338 376961
rect 482282 376887 482338 376896
rect 482204 373966 482324 373994
rect 482296 339697 482324 373966
rect 482388 367577 482416 536794
rect 482468 524476 482520 524482
rect 482468 524418 482520 524424
rect 482374 367568 482430 367577
rect 482374 367503 482430 367512
rect 482376 364404 482428 364410
rect 482376 364346 482428 364352
rect 482282 339688 482338 339697
rect 482282 339623 482338 339632
rect 482388 334937 482416 364346
rect 482480 362953 482508 524418
rect 482560 484424 482612 484430
rect 482560 484366 482612 484372
rect 482466 362944 482522 362953
rect 482466 362879 482522 362888
rect 482572 358329 482600 484366
rect 482652 470620 482704 470626
rect 482652 470562 482704 470568
rect 482558 358320 482614 358329
rect 482558 358255 482614 358264
rect 482664 353705 482692 470562
rect 482744 430636 482796 430642
rect 482744 430578 482796 430584
rect 482650 353696 482706 353705
rect 482650 353631 482706 353640
rect 482756 348945 482784 430578
rect 482836 418192 482888 418198
rect 482836 418134 482888 418140
rect 482742 348936 482798 348945
rect 482742 348871 482798 348880
rect 482848 344321 482876 418134
rect 492692 402286 492720 575878
rect 495084 572354 495112 575892
rect 496740 572422 496768 575892
rect 498396 572762 498424 575892
rect 499592 575878 499974 575906
rect 500972 575878 501630 575906
rect 502352 575878 503286 575906
rect 503732 575878 504942 575906
rect 497464 572756 497516 572762
rect 497464 572698 497516 572704
rect 498384 572756 498436 572762
rect 498384 572698 498436 572704
rect 496728 572416 496780 572422
rect 496728 572358 496780 572364
rect 495072 572348 495124 572354
rect 495072 572290 495124 572296
rect 497476 402354 497504 572698
rect 499592 402422 499620 575878
rect 500972 402490 501000 575878
rect 502352 403646 502380 575878
rect 503732 403714 503760 575878
rect 503720 403708 503772 403714
rect 503720 403650 503772 403656
rect 502340 403640 502392 403646
rect 502340 403582 502392 403588
rect 506492 402558 506520 575892
rect 508148 573782 508176 575892
rect 509804 573850 509832 575892
rect 509792 573844 509844 573850
rect 509792 573786 509844 573792
rect 508136 573776 508188 573782
rect 508136 573718 508188 573724
rect 511460 573646 511488 575892
rect 511448 573640 511500 573646
rect 511448 573582 511500 573588
rect 513116 573510 513144 575892
rect 514680 573714 514708 575892
rect 514668 573708 514720 573714
rect 514668 573650 514720 573656
rect 516336 573578 516364 575892
rect 516324 573572 516376 573578
rect 516324 573514 516376 573520
rect 513104 573504 513156 573510
rect 513104 573446 513156 573452
rect 517992 573442 518020 575892
rect 519648 574054 519676 575892
rect 519636 574048 519688 574054
rect 519636 573990 519688 573996
rect 517980 573436 518032 573442
rect 517980 573378 518032 573384
rect 521304 573306 521332 575892
rect 522868 573374 522896 575892
rect 522856 573368 522908 573374
rect 522856 573310 522908 573316
rect 521292 573300 521344 573306
rect 521292 573242 521344 573248
rect 524524 573238 524552 575892
rect 524512 573232 524564 573238
rect 524512 573174 524564 573180
rect 526180 573170 526208 575892
rect 526168 573164 526220 573170
rect 526168 573106 526220 573112
rect 527836 573102 527864 575892
rect 527824 573096 527876 573102
rect 527824 573038 527876 573044
rect 506480 402552 506532 402558
rect 506480 402494 506532 402500
rect 500960 402484 501012 402490
rect 500960 402426 501012 402432
rect 499580 402416 499632 402422
rect 499580 402358 499632 402364
rect 497464 402348 497516 402354
rect 497464 402290 497516 402296
rect 492680 402280 492732 402286
rect 492680 402222 492732 402228
rect 482928 396024 482980 396030
rect 482928 395966 482980 395972
rect 482940 395593 482968 395966
rect 482926 395584 482982 395593
rect 482926 395519 482982 395528
rect 529216 391950 529244 683130
rect 530596 400926 530624 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 536104 696992 536156 696998
rect 536104 696934 536156 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 533344 643136 533396 643142
rect 533344 643078 533396 643084
rect 530584 400920 530636 400926
rect 530584 400862 530636 400868
rect 482928 391944 482980 391950
rect 482928 391886 482980 391892
rect 529204 391944 529256 391950
rect 529204 391886 529256 391892
rect 482940 390969 482968 391886
rect 482926 390960 482982 390969
rect 482926 390895 482982 390904
rect 533356 386374 533384 643078
rect 536116 396030 536144 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 538864 630692 538916 630698
rect 538864 630634 538916 630640
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 537484 576904 537536 576910
rect 537484 576846 537536 576852
rect 536104 396024 536156 396030
rect 536104 395966 536156 395972
rect 482928 386368 482980 386374
rect 482926 386336 482928 386345
rect 533344 386368 533396 386374
rect 482980 386336 482982 386345
rect 533344 386310 533396 386316
rect 482926 386271 482982 386280
rect 537496 372570 537524 576846
rect 538876 382226 538904 630634
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 538864 382220 538916 382226
rect 538864 382162 538916 382168
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580276 378146 580304 590951
rect 580264 378140 580316 378146
rect 580264 378082 580316 378088
rect 482928 372564 482980 372570
rect 482928 372506 482980 372512
rect 537484 372564 537536 372570
rect 537484 372506 537536 372512
rect 482940 372337 482968 372506
rect 482926 372328 482982 372337
rect 482926 372263 482982 372272
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 482834 344312 482890 344321
rect 482834 344247 482890 344256
rect 482374 334928 482430 334937
rect 482374 334863 482430 334872
rect 482282 330304 482338 330313
rect 482282 330239 482338 330248
rect 482296 325650 482324 330239
rect 482374 325680 482430 325689
rect 482284 325644 482336 325650
rect 482374 325615 482430 325624
rect 580172 325644 580224 325650
rect 482284 325586 482336 325592
rect 482282 320920 482338 320929
rect 482282 320855 482338 320864
rect 482006 316296 482062 316305
rect 482006 316231 482062 316240
rect 481914 265024 481970 265033
rect 481914 264959 481916 264968
rect 481968 264959 481970 264968
rect 481916 264930 481968 264936
rect 482020 259418 482048 316231
rect 482098 311672 482154 311681
rect 482098 311607 482154 311616
rect 482008 259412 482060 259418
rect 482008 259354 482060 259360
rect 340328 258256 340380 258262
rect 340380 258204 340676 258210
rect 340328 258198 340676 258204
rect 340340 258182 340676 258198
rect 341628 258046 341964 258074
rect 342272 258046 343252 258074
rect 344296 258046 344632 258074
rect 345920 258046 345980 258074
rect 340236 256284 340288 256290
rect 340236 256226 340288 256232
rect 340144 255944 340196 255950
rect 340144 255886 340196 255892
rect 339408 255808 339460 255814
rect 339408 255750 339460 255756
rect 338856 255400 338908 255406
rect 338856 255342 338908 255348
rect 337108 253224 337160 253230
rect 337108 253166 337160 253172
rect 337016 201340 337068 201346
rect 337016 201282 337068 201288
rect 338868 3398 338896 255342
rect 340156 9110 340184 255886
rect 340248 13258 340276 256226
rect 341628 255814 341656 258046
rect 340880 255808 340932 255814
rect 340880 255750 340932 255756
rect 341616 255808 341668 255814
rect 341616 255750 341668 255756
rect 340236 13252 340288 13258
rect 340236 13194 340288 13200
rect 340892 10470 340920 255750
rect 342272 11762 342300 258046
rect 344296 255950 344324 258046
rect 345952 256630 345980 258046
rect 346872 258046 347208 258074
rect 348252 258046 348588 258074
rect 349172 258046 349876 258074
rect 350828 258046 351164 258074
rect 351932 258046 352544 258074
rect 353312 258046 353832 258074
rect 354692 258046 355120 258074
rect 356072 258046 356500 258074
rect 357452 258046 357788 258074
rect 358832 258046 359168 258074
rect 360212 258046 360456 258074
rect 361592 258046 361744 258074
rect 362972 258046 363124 258074
rect 345940 256624 345992 256630
rect 345940 256566 345992 256572
rect 344284 255944 344336 255950
rect 344284 255886 344336 255892
rect 345664 255536 345716 255542
rect 345664 255478 345716 255484
rect 342260 11756 342312 11762
rect 342260 11698 342312 11704
rect 340880 10464 340932 10470
rect 340880 10406 340932 10412
rect 340144 9104 340196 9110
rect 340144 9046 340196 9052
rect 345676 9042 345704 255478
rect 346872 255406 346900 258046
rect 347044 256624 347096 256630
rect 347044 256566 347096 256572
rect 346860 255400 346912 255406
rect 346860 255342 346912 255348
rect 347056 202230 347084 256566
rect 348252 255542 348280 258046
rect 348240 255536 348292 255542
rect 348240 255478 348292 255484
rect 347044 202224 347096 202230
rect 347044 202166 347096 202172
rect 349172 10538 349200 258046
rect 350828 256358 350856 258046
rect 350816 256352 350868 256358
rect 350816 256294 350868 256300
rect 349160 10532 349212 10538
rect 349160 10474 349212 10480
rect 345664 9036 345716 9042
rect 345664 8978 345716 8984
rect 351932 4146 351960 258046
rect 352564 256352 352616 256358
rect 352564 256294 352616 256300
rect 352576 200705 352604 256294
rect 352562 200696 352618 200705
rect 352562 200631 352618 200640
rect 353312 4350 353340 258046
rect 354692 5642 354720 258046
rect 354680 5636 354732 5642
rect 354680 5578 354732 5584
rect 353300 4344 353352 4350
rect 353300 4286 353352 4292
rect 351920 4140 351972 4146
rect 351920 4082 351972 4088
rect 356072 3942 356100 258046
rect 357452 4010 357480 258046
rect 358832 4282 358860 258046
rect 360212 13190 360240 258046
rect 361592 256562 361620 258046
rect 361580 256556 361632 256562
rect 361580 256498 361632 256504
rect 360200 13184 360252 13190
rect 360200 13126 360252 13132
rect 362972 7070 363000 258046
rect 364398 257802 364426 258060
rect 365700 258046 365760 258074
rect 367080 258046 367140 258074
rect 364352 257774 364426 257802
rect 362960 7064 363012 7070
rect 362960 7006 363012 7012
rect 364352 4418 364380 257774
rect 365732 256630 365760 258046
rect 365720 256624 365772 256630
rect 365720 256566 365772 256572
rect 367112 256494 367140 258046
rect 367204 258046 368368 258074
rect 369320 258046 369656 258074
rect 369872 258046 371036 258074
rect 371252 258046 372324 258074
rect 373276 258046 373612 258074
rect 374012 258046 374992 258074
rect 375392 258046 376280 258074
rect 376772 258046 377660 258074
rect 378152 258046 378948 258074
rect 379900 258046 380236 258074
rect 380912 258046 381616 258074
rect 382292 258046 382904 258074
rect 383672 258046 384192 258074
rect 385052 258046 385572 258074
rect 386432 258046 386860 258074
rect 387812 258046 388148 258074
rect 389192 258046 389528 258074
rect 390572 258046 390816 258074
rect 391952 258046 392104 258074
rect 393332 258046 393484 258074
rect 367100 256488 367152 256494
rect 367100 256430 367152 256436
rect 364340 4412 364392 4418
rect 364340 4354 364392 4360
rect 358820 4276 358872 4282
rect 358820 4218 358872 4224
rect 367204 4078 367232 258046
rect 369320 256494 369348 258046
rect 367744 256488 367796 256494
rect 367744 256430 367796 256436
rect 369308 256488 369360 256494
rect 369308 256430 369360 256436
rect 367756 203658 367784 256430
rect 367744 203652 367796 203658
rect 367744 203594 367796 203600
rect 369872 51882 369900 258046
rect 370504 255672 370556 255678
rect 370504 255614 370556 255620
rect 370516 203726 370544 255614
rect 370504 203720 370556 203726
rect 370504 203662 370556 203668
rect 369860 51876 369912 51882
rect 369860 51818 369912 51824
rect 367192 4072 367244 4078
rect 367192 4014 367244 4020
rect 357440 4004 357492 4010
rect 357440 3946 357492 3952
rect 356060 3936 356112 3942
rect 356060 3878 356112 3884
rect 371252 3874 371280 258046
rect 373276 255678 373304 258046
rect 373264 255672 373316 255678
rect 373264 255614 373316 255620
rect 374012 51746 374040 258046
rect 374644 256488 374696 256494
rect 374644 256430 374696 256436
rect 374000 51740 374052 51746
rect 374000 51682 374052 51688
rect 374656 9178 374684 256430
rect 374644 9172 374696 9178
rect 374644 9114 374696 9120
rect 371240 3868 371292 3874
rect 371240 3810 371292 3816
rect 375392 3806 375420 258046
rect 376772 29918 376800 258046
rect 376760 29912 376812 29918
rect 376760 29854 376812 29860
rect 378152 13122 378180 258046
rect 379900 256426 379928 258046
rect 379888 256420 379940 256426
rect 379888 256362 379940 256368
rect 380912 29782 380940 258046
rect 382292 51814 382320 258046
rect 382280 51808 382332 51814
rect 382280 51750 382332 51756
rect 380900 29776 380952 29782
rect 380900 29718 380952 29724
rect 378140 13116 378192 13122
rect 378140 13058 378192 13064
rect 383672 7206 383700 258046
rect 385052 29850 385080 258046
rect 385040 29844 385092 29850
rect 385040 29786 385092 29792
rect 383660 7200 383712 7206
rect 383660 7142 383712 7148
rect 386432 7138 386460 258046
rect 387812 7274 387840 258046
rect 389192 8974 389220 258046
rect 390572 256494 390600 258046
rect 390560 256488 390612 256494
rect 390560 256430 390612 256436
rect 389180 8968 389232 8974
rect 389180 8910 389232 8916
rect 387800 7268 387852 7274
rect 387800 7210 387852 7216
rect 386420 7132 386472 7138
rect 386420 7074 386472 7080
rect 375380 3800 375432 3806
rect 375380 3742 375432 3748
rect 391952 3602 391980 258046
rect 393332 29646 393360 258046
rect 394758 257802 394786 258060
rect 396138 257802 396166 258060
rect 397440 258046 397500 258074
rect 394712 257774 394786 257802
rect 396092 257774 396166 257802
rect 393320 29640 393372 29646
rect 393320 29582 393372 29588
rect 394712 5914 394740 257774
rect 396092 7410 396120 257774
rect 397472 256290 397500 258046
rect 397564 258046 398728 258074
rect 398852 258046 400108 258074
rect 400232 258046 401396 258074
rect 401612 258046 402684 258074
rect 402992 258046 404064 258074
rect 405016 258046 405352 258074
rect 405752 258046 406640 258074
rect 407132 258046 408020 258074
rect 408972 258046 409308 258074
rect 409892 258046 410688 258074
rect 411272 258046 411976 258074
rect 412652 258046 413264 258074
rect 414032 258046 414644 258074
rect 415596 258046 415932 258074
rect 416792 258046 417220 258074
rect 418172 258046 418600 258074
rect 419552 258046 419888 258074
rect 420932 258046 421176 258074
rect 422312 258046 422556 258074
rect 423692 258046 423844 258074
rect 397460 256284 397512 256290
rect 397460 256226 397512 256232
rect 396080 7404 396132 7410
rect 396080 7346 396132 7352
rect 394700 5908 394752 5914
rect 394700 5850 394752 5856
rect 397564 5710 397592 258046
rect 397552 5704 397604 5710
rect 397552 5646 397604 5652
rect 398852 3670 398880 258046
rect 400232 29714 400260 258046
rect 400220 29708 400272 29714
rect 400220 29650 400272 29656
rect 401612 5778 401640 258046
rect 402992 7342 403020 258046
rect 405016 256222 405044 258046
rect 405004 256216 405056 256222
rect 405004 256158 405056 256164
rect 402980 7336 403032 7342
rect 402980 7278 403032 7284
rect 405752 5846 405780 258046
rect 407132 7478 407160 258046
rect 408972 256358 409000 258046
rect 408960 256352 409012 256358
rect 408960 256294 409012 256300
rect 407120 7472 407172 7478
rect 407120 7414 407172 7420
rect 409892 6050 409920 258046
rect 411272 7546 411300 258046
rect 412652 10402 412680 258046
rect 412640 10396 412692 10402
rect 412640 10338 412692 10344
rect 411260 7540 411312 7546
rect 411260 7482 411312 7488
rect 409880 6044 409932 6050
rect 409880 5986 409932 5992
rect 414032 5982 414060 258046
rect 415596 256154 415624 258046
rect 415584 256148 415636 256154
rect 415584 256090 415636 256096
rect 414020 5976 414072 5982
rect 414020 5918 414072 5924
rect 405740 5840 405792 5846
rect 405740 5782 405792 5788
rect 401600 5772 401652 5778
rect 401600 5714 401652 5720
rect 416792 4486 416820 258046
rect 418172 6118 418200 258046
rect 419552 8294 419580 258046
rect 419540 8288 419592 8294
rect 419540 8230 419592 8236
rect 418160 6112 418212 6118
rect 418160 6054 418212 6060
rect 420932 4554 420960 258046
rect 422312 6866 422340 258046
rect 423692 8226 423720 258046
rect 425118 257802 425146 258060
rect 426498 257802 426526 258060
rect 427800 258046 427860 258074
rect 429180 258046 429240 258074
rect 425072 257774 425146 257802
rect 426452 257774 426526 257802
rect 423680 8220 423732 8226
rect 423680 8162 423732 8168
rect 422300 6860 422352 6866
rect 422300 6802 422352 6808
rect 425072 4622 425100 257774
rect 426452 6730 426480 257774
rect 427832 8022 427860 258046
rect 427820 8016 427872 8022
rect 427820 7958 427872 7964
rect 426440 6724 426492 6730
rect 426440 6666 426492 6672
rect 429212 5370 429240 258046
rect 429304 258046 430468 258074
rect 430592 258046 431756 258074
rect 431972 258046 433136 258074
rect 433352 258046 434424 258074
rect 434732 258046 435712 258074
rect 436112 258046 437092 258074
rect 437492 258046 438380 258074
rect 438872 258046 439668 258074
rect 440252 258046 441048 258074
rect 441632 258046 442336 258074
rect 443012 258046 443624 258074
rect 444392 258046 445004 258074
rect 445772 258046 446292 258074
rect 447152 258046 447672 258074
rect 448532 258046 448960 258074
rect 449912 258046 450248 258074
rect 451292 258046 451628 258074
rect 452672 258046 452916 258074
rect 454052 258046 454204 258074
rect 455432 258046 455584 258074
rect 429304 6662 429332 258046
rect 430592 8090 430620 258046
rect 430580 8084 430632 8090
rect 430580 8026 430632 8032
rect 429292 6656 429344 6662
rect 429292 6598 429344 6604
rect 429200 5364 429252 5370
rect 429200 5306 429252 5312
rect 431972 4690 432000 258046
rect 433352 6798 433380 258046
rect 434732 8158 434760 258046
rect 434720 8152 434772 8158
rect 434720 8094 434772 8100
rect 433340 6792 433392 6798
rect 433340 6734 433392 6740
rect 436112 5438 436140 258046
rect 436744 256148 436796 256154
rect 436744 256090 436796 256096
rect 436756 202298 436784 256090
rect 436744 202292 436796 202298
rect 436744 202234 436796 202240
rect 437492 6526 437520 258046
rect 437480 6520 437532 6526
rect 437480 6462 437532 6468
rect 436100 5432 436152 5438
rect 436100 5374 436152 5380
rect 431960 4684 432012 4690
rect 431960 4626 432012 4632
rect 425060 4616 425112 4622
rect 425060 4558 425112 4564
rect 420920 4548 420972 4554
rect 420920 4490 420972 4496
rect 416780 4480 416832 4486
rect 416780 4422 416832 4428
rect 398840 3664 398892 3670
rect 398840 3606 398892 3612
rect 391940 3596 391992 3602
rect 391940 3538 391992 3544
rect 438872 3534 438900 258046
rect 440252 5506 440280 258046
rect 441632 6594 441660 258046
rect 443012 7954 443040 258046
rect 443000 7948 443052 7954
rect 443000 7890 443052 7896
rect 441620 6588 441672 6594
rect 441620 6530 441672 6536
rect 440240 5500 440292 5506
rect 440240 5442 440292 5448
rect 444392 4758 444420 258046
rect 445772 6322 445800 258046
rect 445760 6316 445812 6322
rect 445760 6258 445812 6264
rect 444380 4752 444432 4758
rect 444380 4694 444432 4700
rect 438860 3528 438912 3534
rect 438860 3470 438912 3476
rect 447152 3466 447180 258046
rect 448532 5166 448560 258046
rect 449912 6458 449940 258046
rect 451292 7886 451320 258046
rect 451280 7880 451332 7886
rect 451280 7822 451332 7828
rect 449900 6452 449952 6458
rect 449900 6394 449952 6400
rect 452672 5302 452700 258046
rect 454052 6254 454080 258046
rect 455432 256086 455460 258046
rect 456858 257802 456886 258060
rect 458160 258046 458220 258074
rect 459540 258046 459692 258074
rect 456812 257774 456886 257802
rect 455420 256080 455472 256086
rect 455420 256022 455472 256028
rect 454040 6248 454092 6254
rect 454040 6190 454092 6196
rect 452660 5296 452712 5302
rect 452660 5238 452712 5244
rect 448520 5160 448572 5166
rect 448520 5102 448572 5108
rect 456812 4894 456840 257774
rect 458192 203590 458220 258046
rect 459560 253224 459612 253230
rect 459560 253166 459612 253172
rect 458180 203584 458232 203590
rect 458180 203526 458232 203532
rect 459572 5234 459600 253166
rect 459664 7682 459692 258046
rect 460492 258046 460828 258074
rect 460952 258046 462116 258074
rect 463160 258046 463496 258074
rect 463712 258046 464784 258074
rect 465092 258046 466164 258074
rect 466472 258046 467452 258074
rect 467852 258046 468740 258074
rect 469232 258046 470120 258074
rect 470612 258046 471408 258074
rect 471992 258046 472696 258074
rect 473740 258046 474076 258074
rect 475028 258046 475364 258074
rect 476132 258046 476652 258074
rect 477696 258046 478032 258074
rect 478892 258046 479320 258074
rect 460492 253230 460520 258046
rect 460480 253224 460532 253230
rect 460480 253166 460532 253172
rect 459652 7676 459704 7682
rect 459652 7618 459704 7624
rect 460952 6390 460980 258046
rect 463160 256018 463188 258046
rect 463148 256012 463200 256018
rect 463148 255954 463200 255960
rect 460940 6384 460992 6390
rect 460940 6326 460992 6332
rect 459560 5228 459612 5234
rect 459560 5170 459612 5176
rect 463712 4962 463740 258046
rect 465092 202162 465120 258046
rect 465724 256012 465776 256018
rect 465724 255954 465776 255960
rect 465080 202156 465132 202162
rect 465080 202098 465132 202104
rect 463700 4956 463752 4962
rect 463700 4898 463752 4904
rect 456800 4888 456852 4894
rect 456800 4830 456852 4836
rect 465736 3738 465764 255954
rect 466472 7818 466500 258046
rect 466460 7812 466512 7818
rect 466460 7754 466512 7760
rect 467852 5030 467880 258046
rect 469232 6186 469260 258046
rect 470612 7750 470640 258046
rect 470600 7744 470652 7750
rect 470600 7686 470652 7692
rect 469220 6180 469272 6186
rect 469220 6122 469272 6128
rect 471992 5098 472020 258046
rect 473740 256154 473768 258046
rect 473728 256148 473780 256154
rect 473728 256090 473780 256096
rect 475028 256018 475056 258046
rect 475384 256352 475436 256358
rect 475384 256294 475436 256300
rect 475016 256012 475068 256018
rect 475016 255954 475068 255960
rect 475396 10334 475424 256294
rect 475384 10328 475436 10334
rect 475384 10270 475436 10276
rect 471980 5092 472032 5098
rect 471980 5034 472032 5040
rect 467840 5024 467892 5030
rect 467840 4966 467892 4972
rect 476132 4826 476160 258046
rect 477696 256358 477724 258046
rect 477684 256352 477736 256358
rect 477684 256294 477736 256300
rect 478892 7614 478920 258046
rect 482112 233238 482140 311607
rect 482190 307048 482246 307057
rect 482190 306983 482246 306992
rect 482100 233232 482152 233238
rect 482100 233174 482152 233180
rect 482204 219434 482232 306983
rect 482296 273222 482324 320855
rect 482388 313274 482416 325615
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 482376 313268 482428 313274
rect 482376 313210 482428 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 482926 302288 482982 302297
rect 482926 302223 482982 302232
rect 482834 297664 482890 297673
rect 482834 297599 482890 297608
rect 482742 293040 482798 293049
rect 482742 292975 482798 292984
rect 482650 288280 482706 288289
rect 482650 288215 482706 288224
rect 482558 283656 482614 283665
rect 482558 283591 482614 283600
rect 482466 279032 482522 279041
rect 482466 278967 482522 278976
rect 482374 274272 482430 274281
rect 482374 274207 482430 274216
rect 482388 273834 482416 274207
rect 482376 273828 482428 273834
rect 482376 273770 482428 273776
rect 482284 273216 482336 273222
rect 482284 273158 482336 273164
rect 482374 269648 482430 269657
rect 482374 269583 482430 269592
rect 482282 260400 482338 260409
rect 482282 260335 482338 260344
rect 482192 219428 482244 219434
rect 482192 219370 482244 219376
rect 482296 20670 482324 260335
rect 482388 60722 482416 269583
rect 482480 100706 482508 278967
rect 482572 113150 482600 283591
rect 482664 139398 482692 288215
rect 482756 153202 482784 292975
rect 482848 179382 482876 297599
rect 482940 193186 482968 302223
rect 485044 273828 485096 273834
rect 485044 273770 485096 273776
rect 483664 264988 483716 264994
rect 483664 264930 483716 264936
rect 482928 193180 482980 193186
rect 482928 193122 482980 193128
rect 482836 179376 482888 179382
rect 482836 179318 482888 179324
rect 482744 153196 482796 153202
rect 482744 153138 482796 153144
rect 482652 139392 482704 139398
rect 482652 139334 482704 139340
rect 482560 113144 482612 113150
rect 482560 113086 482612 113092
rect 482468 100700 482520 100706
rect 482468 100642 482520 100648
rect 482376 60716 482428 60722
rect 482376 60658 482428 60664
rect 483676 33114 483704 264930
rect 485056 73166 485084 273770
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 485044 73160 485096 73166
rect 485044 73102 485096 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 483664 33108 483716 33114
rect 580170 33079 580172 33088
rect 483664 33050 483716 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 482284 20664 482336 20670
rect 482284 20606 482336 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 478880 7608 478932 7614
rect 478880 7550 478932 7556
rect 476120 4820 476172 4826
rect 476120 4762 476172 4768
rect 465724 3732 465776 3738
rect 465724 3674 465776 3680
rect 447140 3460 447192 3466
rect 447140 3402 447192 3408
rect 338856 3392 338908 3398
rect 338856 3334 338908 3340
rect 336096 3324 336148 3330
rect 336096 3266 336148 3272
rect 334624 3120 334676 3126
rect 334624 3062 334676 3068
rect 324964 2916 325016 2922
rect 324964 2858 325016 2864
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 354 7738 480
rect 8128 462 8206 490
rect 8128 354 8156 462
rect 8772 480 8800 711
rect 9600 649 9628 1158
rect 10980 1057 11008 1226
rect 11704 1148 11756 1154
rect 11704 1090 11756 1096
rect 10966 1048 11022 1057
rect 10966 983 11022 992
rect 11716 921 11744 1090
rect 12346 1048 12402 1057
rect 12346 983 12402 992
rect 11702 912 11758 921
rect 9956 876 10008 882
rect 11702 847 11758 856
rect 9956 818 10008 824
rect 9586 640 9642 649
rect 9586 575 9642 584
rect 9968 480 9996 818
rect 11150 640 11206 649
rect 11150 575 11206 584
rect 11164 480 11192 575
rect 12360 480 12388 983
rect 17052 480 17080 2751
rect 19248 1080 19300 1086
rect 19246 1048 19248 1057
rect 19300 1048 19302 1057
rect 17868 1012 17920 1018
rect 19246 983 19302 992
rect 17868 954 17920 960
rect 17880 785 17908 954
rect 19430 912 19486 921
rect 19430 847 19486 856
rect 17866 776 17922 785
rect 17866 711 17922 720
rect 18234 776 18290 785
rect 18234 711 18290 720
rect 18248 480 18276 711
rect 19444 480 19472 847
rect 8206 439 8262 448
rect 7626 326 8156 354
rect 7626 -960 7738 326
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 82 13626 480
rect 14710 218 14822 480
rect 14568 202 14822 218
rect 14556 196 14822 202
rect 14608 190 14822 196
rect 14556 138 14608 144
rect 13728 128 13780 134
rect 13514 76 13728 82
rect 13514 70 13780 76
rect 13514 54 13768 70
rect 13514 -960 13626 54
rect 14710 -960 14822 190
rect 15906 218 16018 480
rect 16212 264 16264 270
rect 15906 212 16212 218
rect 15906 206 16264 212
rect 15906 190 16252 206
rect 15906 -960 16018 190
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20364 105 20392 2774
rect 20598 354 20710 480
rect 20456 338 20710 354
rect 20444 332 20710 338
rect 20496 326 20710 332
rect 20444 274 20496 280
rect 20350 96 20406 105
rect 20350 31 20406 40
rect 20598 -960 20710 326
rect 21468 241 21496 2774
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 21836 480 21864 983
rect 21454 232 21510 241
rect 21454 167 21510 176
rect 21794 -960 21906 480
rect 22572 377 22600 2774
rect 23722 2802 23750 3060
rect 24826 2802 24854 3060
rect 25930 2802 25958 3060
rect 27034 2802 27062 3060
rect 28138 2802 28166 3060
rect 29242 2802 29270 3060
rect 23018 2751 23074 2760
rect 23676 2774 23750 2802
rect 24780 2774 24854 2802
rect 25884 2774 25958 2802
rect 26988 2774 27062 2802
rect 28092 2774 28166 2802
rect 29196 2774 29270 2802
rect 30104 2848 30156 2854
rect 30346 2802 30374 3060
rect 31450 2802 31478 3060
rect 30104 2790 30156 2796
rect 23032 480 23060 2751
rect 23676 1222 23704 2774
rect 23664 1216 23716 1222
rect 23664 1158 23716 1164
rect 23848 1216 23900 1222
rect 23848 1158 23900 1164
rect 23860 1057 23888 1158
rect 24780 1154 24808 2774
rect 25884 1290 25912 2774
rect 25872 1284 25924 1290
rect 25872 1226 25924 1232
rect 24768 1148 24820 1154
rect 24768 1090 24820 1096
rect 23846 1048 23902 1057
rect 23846 983 23902 992
rect 25780 944 25832 950
rect 25780 886 25832 892
rect 22558 368 22614 377
rect 22558 303 22614 312
rect 22990 -960 23102 480
rect 24186 354 24298 480
rect 24766 368 24822 377
rect 24186 326 24766 354
rect 24186 -960 24298 326
rect 24766 303 24822 312
rect 25290 354 25402 480
rect 25792 354 25820 886
rect 26988 513 27016 2774
rect 28092 1018 28120 2774
rect 28264 1352 28316 1358
rect 28264 1294 28316 1300
rect 28080 1012 28132 1018
rect 28080 954 28132 960
rect 28276 649 28304 1294
rect 29196 882 29224 2774
rect 29184 876 29236 882
rect 29184 818 29236 824
rect 28262 640 28318 649
rect 28262 575 28318 584
rect 26974 504 27030 513
rect 25290 326 25820 354
rect 25290 -960 25402 326
rect 26330 232 26386 241
rect 26486 218 26598 480
rect 28170 504 28226 513
rect 26974 439 27030 448
rect 26386 190 26598 218
rect 26330 167 26386 176
rect 26486 -960 26598 190
rect 27682 354 27794 480
rect 30116 480 30144 2790
rect 30300 2774 30374 2802
rect 31404 2774 31478 2802
rect 32554 2802 32582 3060
rect 33658 2802 33686 3060
rect 34762 2802 34790 3060
rect 35866 2961 35894 3060
rect 35852 2952 35908 2961
rect 35852 2887 35908 2896
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 32554 2774 32628 2802
rect 30300 1358 30328 2774
rect 30288 1352 30340 1358
rect 30288 1294 30340 1300
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 30288 1148 30340 1154
rect 30288 1090 30340 1096
rect 28170 439 28226 448
rect 28184 354 28212 439
rect 27682 326 28212 354
rect 28724 400 28776 406
rect 28878 354 28990 480
rect 28776 348 28990 354
rect 28724 342 28990 348
rect 28736 326 28990 342
rect 27682 -960 27794 326
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30300 377 30328 1090
rect 31036 921 31064 1294
rect 31404 1086 31432 2774
rect 31392 1080 31444 1086
rect 31392 1022 31444 1028
rect 31022 912 31078 921
rect 31022 847 31078 856
rect 31298 640 31354 649
rect 31298 575 31354 584
rect 31312 480 31340 575
rect 30286 368 30342 377
rect 30286 303 30342 312
rect 31270 -960 31382 480
rect 32220 468 32272 474
rect 32220 410 32272 416
rect 32232 354 32260 410
rect 32374 354 32486 480
rect 32232 326 32486 354
rect 32374 -960 32486 326
rect 32600 134 32628 2774
rect 33428 2774 33686 2802
rect 34624 2774 34790 2802
rect 33232 1012 33284 1018
rect 33232 954 33284 960
rect 33244 649 33272 954
rect 33230 640 33286 649
rect 33230 575 33286 584
rect 33428 202 33456 2774
rect 33612 598 33824 626
rect 33612 480 33640 598
rect 33416 196 33468 202
rect 33416 138 33468 144
rect 32588 128 32640 134
rect 32588 70 32640 76
rect 33570 -960 33682 480
rect 33796 134 33824 598
rect 34624 270 34652 2774
rect 34794 2544 34850 2553
rect 34794 2479 34850 2488
rect 34808 480 34836 2479
rect 36004 480 36032 2858
rect 36970 2802 36998 3060
rect 36924 2774 36998 2802
rect 37188 2848 37240 2854
rect 38074 2802 38102 3060
rect 39178 2802 39206 3060
rect 40282 2802 40310 3060
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 37188 2790 37240 2796
rect 36924 785 36952 2774
rect 37200 1290 37228 2790
rect 38028 2774 38102 2802
rect 39132 2774 39206 2802
rect 40236 2774 40310 2802
rect 38028 1358 38056 2774
rect 38016 1352 38068 1358
rect 38016 1294 38068 1300
rect 37188 1284 37240 1290
rect 37188 1226 37240 1232
rect 37004 1080 37056 1086
rect 37004 1022 37056 1028
rect 36910 776 36966 785
rect 36910 711 36966 720
rect 37016 513 37044 1022
rect 37002 504 37058 513
rect 34612 264 34664 270
rect 34612 206 34664 212
rect 33784 128 33836 134
rect 33784 70 33836 76
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37002 439 37058 448
rect 37158 218 37270 480
rect 37016 202 37270 218
rect 37004 196 37270 202
rect 37056 190 37270 196
rect 37004 138 37056 144
rect 37158 -960 37270 190
rect 38354 218 38466 480
rect 39132 338 39160 2774
rect 40236 1222 40264 2774
rect 40420 1222 40448 2858
rect 41386 2825 41414 3060
rect 41880 2848 41932 2854
rect 41372 2816 41428 2825
rect 42490 2802 42518 3060
rect 43594 2802 43622 3060
rect 44698 2802 44726 3060
rect 45802 2802 45830 3060
rect 46906 2802 46934 3060
rect 48010 2802 48038 3060
rect 49114 2802 49142 3060
rect 41880 2790 41932 2796
rect 41372 2751 41428 2760
rect 40774 2680 40830 2689
rect 40696 2638 40774 2666
rect 40224 1216 40276 1222
rect 40224 1158 40276 1164
rect 40408 1216 40460 1222
rect 40408 1158 40460 1164
rect 40696 480 40724 2638
rect 40774 2615 40830 2624
rect 41892 480 41920 2790
rect 42444 2774 42518 2802
rect 43548 2774 43622 2802
rect 44652 2774 44726 2802
rect 45756 2774 45830 2802
rect 46860 2774 46934 2802
rect 47964 2774 48038 2802
rect 49068 2774 49142 2802
rect 49608 2848 49660 2854
rect 50218 2802 50246 3060
rect 51322 2938 51350 3060
rect 52426 2961 52454 3060
rect 49608 2790 49660 2796
rect 42444 1154 42472 2774
rect 42432 1148 42484 1154
rect 42432 1090 42484 1096
rect 43548 950 43576 2774
rect 43536 944 43588 950
rect 43536 886 43588 892
rect 42892 536 42944 542
rect 39550 354 39662 480
rect 39408 338 39662 354
rect 39120 332 39172 338
rect 39120 274 39172 280
rect 39396 332 39662 338
rect 39448 326 39662 332
rect 39396 274 39448 280
rect 38568 264 38620 270
rect 38354 212 38568 218
rect 38354 206 38620 212
rect 38354 190 38608 206
rect 38354 -960 38466 190
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42892 478 42944 484
rect 42904 354 42932 478
rect 43046 354 43158 480
rect 42904 326 43158 354
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 44652 241 44680 2774
rect 45756 1086 45784 2774
rect 45744 1080 45796 1086
rect 45744 1022 45796 1028
rect 46664 672 46716 678
rect 46664 614 46716 620
rect 45468 604 45520 610
rect 45468 546 45520 552
rect 45480 480 45508 546
rect 46676 480 46704 614
rect 44638 232 44694 241
rect 44638 167 44694 176
rect 44638 96 44694 105
rect 44242 54 44638 82
rect 44242 -960 44354 54
rect 44638 31 44694 40
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 46860 406 46888 2774
rect 47858 2680 47914 2689
rect 47858 2615 47914 2624
rect 47872 480 47900 2615
rect 47964 1290 47992 2774
rect 47952 1284 48004 1290
rect 47952 1226 48004 1232
rect 49068 1018 49096 2774
rect 49620 1290 49648 2790
rect 49988 2774 50246 2802
rect 51184 2910 51350 2938
rect 52412 2952 52468 2961
rect 49608 1284 49660 1290
rect 49608 1226 49660 1232
rect 49056 1012 49108 1018
rect 49056 954 49108 960
rect 46848 400 46900 406
rect 46848 342 46900 348
rect 47830 -960 47942 480
rect 48780 400 48832 406
rect 48934 354 49046 480
rect 49988 474 50016 2774
rect 50160 740 50212 746
rect 50160 682 50212 688
rect 50172 480 50200 682
rect 49976 468 50028 474
rect 49976 410 50028 416
rect 48832 348 49046 354
rect 48780 342 49046 348
rect 48792 326 49046 342
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51184 134 51212 2910
rect 52412 2887 52468 2896
rect 51356 2848 51408 2854
rect 53530 2802 53558 3060
rect 54634 2802 54662 3060
rect 55738 2802 55766 3060
rect 56842 2802 56870 3060
rect 57946 2825 57974 3060
rect 51356 2790 51408 2796
rect 51368 480 51396 2790
rect 53484 2774 53558 2802
rect 54588 2774 54662 2802
rect 55692 2774 55766 2802
rect 56796 2774 56870 2802
rect 57932 2816 57988 2825
rect 53010 2680 53066 2689
rect 53010 2615 53066 2624
rect 51172 128 51224 134
rect 51172 70 51224 76
rect 51326 -960 51438 480
rect 52522 354 52634 480
rect 53024 354 53052 2615
rect 53484 1222 53512 2774
rect 53472 1216 53524 1222
rect 53472 1158 53524 1164
rect 52522 326 53052 354
rect 52522 -960 52634 326
rect 53564 128 53616 134
rect 53718 82 53830 480
rect 54588 202 54616 2774
rect 54914 218 55026 480
rect 55692 270 55720 2774
rect 55680 264 55732 270
rect 54914 202 55168 218
rect 55680 206 55732 212
rect 56018 218 56130 480
rect 56796 338 56824 2774
rect 57932 2751 57988 2760
rect 58438 2816 58494 2825
rect 59050 2802 59078 3060
rect 58438 2751 58494 2760
rect 59004 2774 59078 2802
rect 59268 2848 59320 2854
rect 60154 2802 60182 3060
rect 59268 2790 59320 2796
rect 58452 480 58480 2751
rect 59004 1290 59032 2774
rect 59280 1358 59308 2790
rect 60108 2774 60182 2802
rect 60832 2848 60884 2854
rect 61258 2802 61286 3060
rect 62362 2802 62390 3060
rect 63466 2802 63494 3060
rect 60832 2790 60884 2796
rect 59634 2000 59690 2009
rect 59634 1935 59690 1944
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 58992 1284 59044 1290
rect 58992 1226 59044 1232
rect 59648 480 59676 1935
rect 60108 542 60136 2774
rect 60096 536 60148 542
rect 57214 354 57326 480
rect 57072 338 57326 354
rect 56784 332 56836 338
rect 56784 274 56836 280
rect 57060 332 57326 338
rect 57112 326 57326 332
rect 57060 274 57112 280
rect 56416 264 56468 270
rect 56018 212 56416 218
rect 56018 206 56468 212
rect 54576 196 54628 202
rect 54576 138 54628 144
rect 54914 196 55180 202
rect 54914 190 55128 196
rect 53616 76 53830 82
rect 53564 70 53830 76
rect 53576 54 53830 70
rect 53718 -960 53830 54
rect 54914 -960 55026 190
rect 55128 138 55180 144
rect 56018 190 56456 206
rect 56018 -960 56130 190
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60096 478 60148 484
rect 60844 480 60872 2790
rect 61212 2774 61286 2802
rect 62316 2774 62390 2802
rect 63420 2774 63494 2802
rect 64326 2816 64382 2825
rect 60802 -960 60914 480
rect 61212 105 61240 2774
rect 62316 610 62344 2774
rect 63420 678 63448 2774
rect 64570 2802 64598 3060
rect 64382 2774 64598 2802
rect 65674 2802 65702 3060
rect 66778 2802 66806 3060
rect 67882 2802 67910 3060
rect 68986 2961 69014 3060
rect 68972 2952 69028 2961
rect 68972 2887 69028 2896
rect 65674 2774 65748 2802
rect 64326 2751 64382 2760
rect 65522 2136 65578 2145
rect 65522 2071 65578 2080
rect 63408 672 63460 678
rect 63408 614 63460 620
rect 62304 604 62356 610
rect 62304 546 62356 552
rect 64328 604 64380 610
rect 64328 546 64380 552
rect 63408 536 63460 542
rect 61844 468 61896 474
rect 61844 410 61896 416
rect 61856 354 61884 410
rect 61998 354 62110 480
rect 61856 326 62110 354
rect 61198 96 61254 105
rect 61198 31 61254 40
rect 61998 -960 62110 326
rect 63194 354 63306 480
rect 63408 478 63460 484
rect 64340 480 64368 546
rect 65536 480 65564 2071
rect 63420 354 63448 478
rect 63194 326 63448 354
rect 63194 -960 63306 326
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 65720 406 65748 2774
rect 66732 2774 66806 2802
rect 67836 2774 67910 2802
rect 68928 2848 68980 2854
rect 70090 2802 70118 3060
rect 68928 2790 68980 2796
rect 66732 746 66760 2774
rect 66994 2272 67050 2281
rect 66824 2230 66994 2258
rect 66720 740 66772 746
rect 66720 682 66772 688
rect 66824 626 66852 2230
rect 66994 2207 67050 2216
rect 67836 1358 67864 2774
rect 68940 1358 68968 2790
rect 70044 2774 70118 2802
rect 70308 2848 70360 2854
rect 71194 2802 71222 3060
rect 72298 2802 72326 3060
rect 73402 2802 73430 3060
rect 74506 2961 74534 3060
rect 74492 2952 74548 2961
rect 74492 2887 74548 2896
rect 75610 2802 75638 3060
rect 70308 2790 70360 2796
rect 69110 2408 69166 2417
rect 69110 2343 69166 2352
rect 67824 1352 67876 1358
rect 67824 1294 67876 1300
rect 68928 1352 68980 1358
rect 68928 1294 68980 1300
rect 67916 1216 67968 1222
rect 67916 1158 67968 1164
rect 66732 598 66852 626
rect 66732 480 66760 598
rect 67928 480 67956 1158
rect 69124 480 69152 2343
rect 65708 400 65760 406
rect 65708 342 65760 348
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70044 134 70072 2774
rect 70320 480 70348 2790
rect 71148 2774 71222 2802
rect 72252 2774 72326 2802
rect 73356 2774 73430 2802
rect 75564 2774 75638 2802
rect 76194 2816 76250 2825
rect 70032 128 70084 134
rect 70032 70 70084 76
rect 70278 -960 70390 480
rect 71148 202 71176 2774
rect 71136 196 71188 202
rect 71136 138 71188 144
rect 71474 82 71586 480
rect 72252 270 72280 2774
rect 72606 2544 72662 2553
rect 72606 2479 72662 2488
rect 72620 480 72648 2479
rect 72240 264 72292 270
rect 72240 206 72292 212
rect 71688 128 71740 134
rect 71474 76 71688 82
rect 71474 70 71740 76
rect 71474 54 71728 70
rect 71474 -960 71586 54
rect 72578 -960 72690 480
rect 73356 338 73384 2774
rect 75564 2009 75592 2774
rect 76714 2802 76742 3060
rect 76194 2751 76250 2760
rect 76668 2774 76742 2802
rect 77208 2848 77260 2854
rect 77818 2802 77846 3060
rect 78922 2802 78950 3060
rect 80026 2802 80054 3060
rect 81130 2802 81158 3060
rect 77208 2790 77260 2796
rect 75550 2000 75606 2009
rect 75550 1935 75606 1944
rect 76208 480 76236 2751
rect 76668 1358 76696 2774
rect 76656 1352 76708 1358
rect 76656 1294 76708 1300
rect 77220 1290 77248 2790
rect 77772 2774 77846 2802
rect 78876 2774 78950 2802
rect 79980 2774 80054 2802
rect 81084 2774 81158 2802
rect 82084 2848 82136 2854
rect 82234 2802 82262 3060
rect 83338 2802 83366 3060
rect 84442 2802 84470 3060
rect 85546 2802 85574 3060
rect 86650 2802 86678 3060
rect 87754 2802 87782 3060
rect 88858 2802 88886 3060
rect 89962 2802 89990 3060
rect 91066 2825 91094 3060
rect 82084 2790 82136 2796
rect 77208 1284 77260 1290
rect 77208 1226 77260 1232
rect 77390 640 77446 649
rect 77390 575 77446 584
rect 77404 480 77432 575
rect 73344 332 73396 338
rect 73344 274 73396 280
rect 73774 218 73886 480
rect 73632 202 73886 218
rect 73620 196 73886 202
rect 73672 190 73886 196
rect 73620 138 73672 144
rect 73774 -960 73886 190
rect 74970 218 75082 480
rect 75368 264 75420 270
rect 74970 212 75368 218
rect 74970 206 75420 212
rect 74970 190 75408 206
rect 74970 -960 75082 190
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 77772 474 77800 2774
rect 78876 542 78904 2774
rect 79980 610 80008 2774
rect 81084 2145 81112 2774
rect 81070 2136 81126 2145
rect 81070 2071 81126 2080
rect 81440 1216 81492 1222
rect 81440 1158 81492 1164
rect 79968 604 80020 610
rect 79968 546 80020 552
rect 78864 536 78916 542
rect 77760 468 77812 474
rect 77760 410 77812 416
rect 78404 400 78456 406
rect 78558 354 78670 480
rect 78864 478 78916 484
rect 79662 354 79774 480
rect 78456 348 78670 354
rect 78404 342 78670 348
rect 78416 326 78670 342
rect 79520 338 79774 354
rect 78558 -960 78670 326
rect 79508 332 79774 338
rect 79560 326 79774 332
rect 79508 274 79560 280
rect 79662 -960 79774 326
rect 80858 354 80970 480
rect 81452 354 81480 1158
rect 82096 480 82124 2790
rect 82188 2774 82262 2802
rect 83292 2774 83366 2802
rect 84396 2774 84470 2802
rect 85500 2774 85574 2802
rect 86604 2774 86678 2802
rect 87708 2774 87782 2802
rect 88812 2774 88886 2802
rect 89916 2774 89990 2802
rect 91052 2816 91108 2825
rect 82188 2281 82216 2774
rect 82174 2272 82230 2281
rect 82174 2207 82230 2216
rect 83292 1358 83320 2774
rect 84396 2417 84424 2774
rect 84382 2408 84438 2417
rect 84382 2343 84438 2352
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 85500 1290 85528 2774
rect 85488 1284 85540 1290
rect 85488 1226 85540 1232
rect 83292 598 83504 626
rect 83292 480 83320 598
rect 83476 513 83504 598
rect 84488 598 84700 626
rect 83462 504 83518 513
rect 80858 326 81480 354
rect 80858 -960 80970 326
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84488 480 84516 598
rect 83462 439 83518 448
rect 84446 -960 84558 480
rect 84672 377 84700 598
rect 84658 368 84714 377
rect 84658 303 84714 312
rect 85642 354 85754 480
rect 86132 468 86184 474
rect 86132 410 86184 416
rect 86144 354 86172 410
rect 85642 326 86172 354
rect 85642 -960 85754 326
rect 86604 134 86632 2774
rect 87708 2553 87736 2774
rect 87694 2544 87750 2553
rect 87694 2479 87750 2488
rect 86592 128 86644 134
rect 86592 70 86644 76
rect 86684 128 86736 134
rect 86838 82 86950 480
rect 87786 368 87842 377
rect 87942 354 88054 480
rect 87842 326 88054 354
rect 87786 303 87842 312
rect 86736 76 86950 82
rect 86684 70 86950 76
rect 86696 54 86950 70
rect 86838 -960 86950 54
rect 87942 -960 88054 326
rect 88812 202 88840 2774
rect 89138 218 89250 480
rect 89916 270 89944 2774
rect 91052 2751 91108 2760
rect 91558 2816 91614 2825
rect 92170 2802 92198 3060
rect 93274 2802 93302 3060
rect 94378 2802 94406 3060
rect 95482 2802 95510 3060
rect 96586 2854 96614 3060
rect 91558 2751 91614 2760
rect 92124 2774 92198 2802
rect 93228 2774 93302 2802
rect 94332 2774 94406 2802
rect 95436 2774 95510 2802
rect 96574 2848 96626 2854
rect 97690 2802 97718 3060
rect 96574 2790 96626 2796
rect 97644 2774 97718 2802
rect 98794 2802 98822 3060
rect 99898 2802 99926 3060
rect 101002 2802 101030 3060
rect 102106 2802 102134 3060
rect 103210 2802 103238 3060
rect 104314 2802 104342 3060
rect 105418 2825 105446 3060
rect 98794 2774 98868 2802
rect 99898 2774 99972 2802
rect 91572 480 91600 2751
rect 92124 649 92152 2774
rect 92110 640 92166 649
rect 92110 575 92166 584
rect 89904 264 89956 270
rect 89138 202 89576 218
rect 89904 206 89956 212
rect 88800 196 88852 202
rect 88800 138 88852 144
rect 89138 196 89588 202
rect 89138 190 89536 196
rect 89138 -960 89250 190
rect 89536 138 89588 144
rect 90178 96 90234 105
rect 90334 82 90446 480
rect 90234 54 90446 82
rect 90178 31 90234 40
rect 90334 -960 90446 54
rect 91530 -960 91642 480
rect 92572 264 92624 270
rect 92726 218 92838 480
rect 93228 406 93256 2774
rect 93950 2000 94006 2009
rect 93950 1935 94006 1944
rect 93964 480 93992 1935
rect 93216 400 93268 406
rect 93216 342 93268 348
rect 92624 212 92838 218
rect 92572 206 92838 212
rect 92584 190 92838 206
rect 92726 -960 92838 190
rect 93922 -960 94034 480
rect 94332 338 94360 2774
rect 95436 1222 95464 2774
rect 95424 1216 95476 1222
rect 95424 1158 95476 1164
rect 97644 513 97672 2774
rect 97908 1216 97960 1222
rect 97908 1158 97960 1164
rect 97630 504 97686 513
rect 95118 354 95230 480
rect 94976 338 95230 354
rect 96068 400 96120 406
rect 96222 354 96334 480
rect 96120 348 96334 354
rect 96068 342 96334 348
rect 94320 332 94372 338
rect 94320 274 94372 280
rect 94964 332 95230 338
rect 95016 326 95230 332
rect 96080 326 96334 342
rect 94964 274 95016 280
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 354 97530 480
rect 97630 439 97686 448
rect 97920 354 97948 1158
rect 98644 672 98696 678
rect 98644 614 98696 620
rect 98656 480 98684 614
rect 98840 513 98868 2774
rect 99746 2272 99802 2281
rect 99746 2207 99802 2216
rect 99760 626 99788 2207
rect 99760 598 99880 626
rect 99944 610 99972 2774
rect 100864 2774 101030 2802
rect 102060 2774 102134 2802
rect 103164 2774 103238 2802
rect 104176 2774 104342 2802
rect 105404 2816 105460 2825
rect 98826 504 98882 513
rect 97418 326 97948 354
rect 97418 -960 97530 326
rect 98614 -960 98726 480
rect 99852 480 99880 598
rect 99932 604 99984 610
rect 99932 546 99984 552
rect 98826 439 98882 448
rect 99810 -960 99922 480
rect 100864 134 100892 2774
rect 101034 2136 101090 2145
rect 101034 2071 101090 2080
rect 101048 480 101076 2071
rect 102060 785 102088 2774
rect 102230 2408 102286 2417
rect 102230 2343 102286 2352
rect 102046 776 102102 785
rect 102046 711 102102 720
rect 102244 480 102272 2343
rect 100852 128 100904 134
rect 100852 70 100904 76
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103164 202 103192 2774
rect 103152 196 103204 202
rect 103152 138 103204 144
rect 103306 82 103418 480
rect 103520 128 103572 134
rect 103306 76 103520 82
rect 104176 105 104204 2774
rect 106522 2802 106550 3060
rect 107626 2802 107654 3060
rect 108730 2802 108758 3060
rect 109834 2802 109862 3060
rect 110938 2802 110966 3060
rect 112042 2802 112070 3060
rect 113146 2802 113174 3060
rect 114250 2802 114278 3060
rect 115354 2802 115382 3060
rect 116458 2802 116486 3060
rect 117562 2802 117590 3060
rect 105404 2751 105460 2760
rect 106476 2774 106550 2802
rect 107580 2774 107654 2802
rect 108684 2774 108758 2802
rect 109788 2774 109862 2802
rect 110892 2774 110966 2802
rect 111996 2774 112070 2802
rect 113100 2774 113174 2802
rect 114204 2774 114278 2802
rect 115308 2774 115382 2802
rect 116228 2774 116486 2802
rect 117516 2774 117590 2802
rect 117686 2816 117742 2825
rect 105726 2544 105782 2553
rect 105726 2479 105782 2488
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 104544 480 104572 1294
rect 105740 480 105768 2479
rect 103306 70 103572 76
rect 104162 96 104218 105
rect 103306 54 103560 70
rect 103306 -960 103418 54
rect 104162 31 104218 40
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 270 106504 2774
rect 107580 2009 107608 2774
rect 107566 2000 107622 2009
rect 107566 1935 107622 1944
rect 108118 2000 108174 2009
rect 108118 1935 108174 1944
rect 107200 1284 107252 1290
rect 107200 1226 107252 1232
rect 107212 626 107240 1226
rect 106936 598 107240 626
rect 106936 480 106964 598
rect 108132 480 108160 1935
rect 106464 264 106516 270
rect 106464 206 106516 212
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 108684 338 108712 2774
rect 109314 2680 109370 2689
rect 109314 2615 109370 2624
rect 109328 480 109356 2615
rect 108672 332 108724 338
rect 108672 274 108724 280
rect 109286 -960 109398 480
rect 109788 406 109816 2774
rect 110892 1222 110920 2774
rect 111614 1864 111670 1873
rect 111614 1799 111670 1808
rect 110880 1216 110932 1222
rect 110880 1158 110932 1164
rect 110972 1148 111024 1154
rect 110972 1090 111024 1096
rect 109776 400 109828 406
rect 109776 342 109828 348
rect 110482 354 110594 480
rect 110984 354 111012 1090
rect 111628 480 111656 1799
rect 111996 678 112024 2774
rect 113100 2281 113128 2774
rect 113086 2272 113142 2281
rect 113086 2207 113142 2216
rect 114204 2145 114232 2774
rect 115308 2417 115336 2774
rect 115294 2408 115350 2417
rect 115294 2343 115350 2352
rect 114190 2136 114246 2145
rect 114190 2071 114246 2080
rect 115202 2136 115258 2145
rect 115202 2071 115258 2080
rect 112810 1728 112866 1737
rect 112810 1663 112866 1672
rect 111984 672 112036 678
rect 111984 614 112036 620
rect 112824 480 112852 1663
rect 115216 480 115244 2071
rect 110482 326 111012 354
rect 110482 -960 110594 326
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 218 114090 480
rect 113978 202 114416 218
rect 113978 196 114428 202
rect 113978 190 114376 196
rect 113978 -960 114090 190
rect 114376 138 114428 144
rect 115174 -960 115286 480
rect 116228 134 116256 2774
rect 117516 1358 117544 2774
rect 118666 2802 118694 3060
rect 119770 2802 119798 3060
rect 120874 2802 120902 3060
rect 121978 2802 122006 3060
rect 123082 2802 123110 3060
rect 124186 2802 124214 3060
rect 125290 2802 125318 3060
rect 126394 2802 126422 3060
rect 127498 2802 127526 3060
rect 128602 2802 128630 3060
rect 129706 2825 129734 3060
rect 117686 2751 117742 2760
rect 118620 2774 118694 2802
rect 119724 2774 119798 2802
rect 120828 2774 120902 2802
rect 121932 2774 122006 2802
rect 123036 2774 123110 2802
rect 124140 2774 124214 2802
rect 125244 2774 125318 2802
rect 126348 2774 126422 2802
rect 127452 2774 127526 2802
rect 128556 2774 128630 2802
rect 129692 2816 129748 2825
rect 117700 1442 117728 2751
rect 118620 2553 118648 2774
rect 118606 2544 118662 2553
rect 118606 2479 118662 2488
rect 117608 1414 117728 1442
rect 117504 1352 117556 1358
rect 117504 1294 117556 1300
rect 116492 1216 116544 1222
rect 116492 1158 116544 1164
rect 116504 626 116532 1158
rect 116412 598 116532 626
rect 116412 480 116440 598
rect 117608 480 117636 1414
rect 119724 1290 119752 2774
rect 120828 2009 120856 2774
rect 121932 2689 121960 2774
rect 121918 2680 121974 2689
rect 121918 2615 121974 2624
rect 120814 2000 120870 2009
rect 120814 1935 120870 1944
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 119712 1284 119764 1290
rect 119712 1226 119764 1232
rect 119908 480 119936 1294
rect 121368 1284 121420 1290
rect 121368 1226 121420 1232
rect 121380 626 121408 1226
rect 123036 1154 123064 2774
rect 124140 1873 124168 2774
rect 124126 1864 124182 1873
rect 124126 1799 124182 1808
rect 125244 1737 125272 2774
rect 125230 1728 125286 1737
rect 125230 1663 125286 1672
rect 123024 1148 123076 1154
rect 123024 1090 123076 1096
rect 125140 1148 125192 1154
rect 125140 1090 125192 1096
rect 123482 776 123538 785
rect 123482 711 123538 720
rect 121104 598 121408 626
rect 121104 480 121132 598
rect 123496 480 123524 711
rect 116216 128 116268 134
rect 116216 70 116268 76
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 82 118874 480
rect 119158 96 119214 105
rect 118762 54 119158 82
rect 118762 -960 118874 54
rect 119158 31 119214 40
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 127176 377 127204 598
rect 129384 480 129412 847
rect 130566 640 130622 649
rect 130566 575 130622 584
rect 130580 480 130608 575
rect 130764 513 130792 2774
rect 131868 1426 131896 2774
rect 131856 1420 131908 1426
rect 131856 1362 131908 1368
rect 132040 1352 132092 1358
rect 132040 1294 132092 1300
rect 132052 762 132080 1294
rect 132972 1290 133000 2774
rect 132960 1284 133012 1290
rect 132960 1226 133012 1232
rect 132774 1048 132830 1057
rect 132774 983 132830 992
rect 131776 734 132080 762
rect 130750 504 130806 513
rect 127162 368 127218 377
rect 127162 303 127218 312
rect 128146 218 128258 480
rect 128146 202 128400 218
rect 128146 196 128412 202
rect 128146 190 128360 196
rect 128146 -960 128258 190
rect 128360 138 128412 144
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131776 480 131804 734
rect 132788 649 132816 983
rect 132774 640 132830 649
rect 132774 575 132830 584
rect 132958 640 133014 649
rect 132958 575 133014 584
rect 132972 480 133000 575
rect 130750 439 130806 448
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133984 134 134012 2774
rect 134352 1442 134380 2858
rect 135226 2802 135254 3060
rect 136330 2802 136358 3060
rect 137434 2802 137462 3060
rect 138538 2802 138566 3060
rect 139642 2802 139670 3060
rect 140746 2802 140774 3060
rect 141850 2802 141878 3060
rect 142954 2802 142982 3060
rect 144058 2802 144086 3060
rect 145162 2922 145190 3060
rect 145150 2916 145202 2922
rect 145150 2858 145202 2864
rect 146266 2802 146294 3060
rect 134168 1414 134380 1442
rect 135180 2774 135254 2802
rect 136284 2774 136358 2802
rect 137296 2774 137462 2802
rect 138492 2774 138566 2802
rect 139596 2774 139670 2802
rect 140700 2774 140774 2802
rect 141804 2774 141878 2802
rect 142908 2774 142982 2802
rect 144012 2774 144086 2802
rect 146220 2774 146294 2802
rect 147126 2816 147182 2825
rect 134168 480 134196 1414
rect 135180 785 135208 2774
rect 135258 2000 135314 2009
rect 135258 1935 135314 1944
rect 135166 776 135222 785
rect 135166 711 135222 720
rect 135272 480 135300 1935
rect 136284 1222 136312 2774
rect 136272 1216 136324 1222
rect 136272 1158 136324 1164
rect 136454 776 136510 785
rect 136454 711 136510 720
rect 136468 480 136496 711
rect 133972 128 134024 134
rect 133972 70 134024 76
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 218 144818 480
rect 144706 202 144960 218
rect 144706 196 144972 202
rect 144706 190 144920 196
rect 144706 -960 144818 190
rect 144920 138 144972 144
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 148506 439 148562 448
rect 149348 134 149376 2774
rect 149518 2544 149574 2553
rect 149518 2479 149574 2488
rect 149532 480 149560 2479
rect 149336 128 149388 134
rect 149336 70 149388 76
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155052 202 155080 2774
rect 155406 2272 155462 2281
rect 155406 2207 155462 2216
rect 155420 480 155448 2207
rect 156156 1358 156184 2774
rect 158410 2802 158438 3060
rect 159514 2802 159542 3060
rect 160618 2802 160646 3060
rect 161722 2802 161750 3060
rect 162826 2854 162854 3060
rect 157292 2751 157348 2760
rect 158364 2774 158438 2802
rect 159468 2774 159542 2802
rect 160572 2774 160646 2802
rect 161676 2774 161750 2802
rect 162814 2848 162866 2854
rect 163930 2802 163958 3060
rect 165034 2802 165062 3060
rect 166138 2802 166166 3060
rect 167242 2802 167270 3060
rect 168346 2802 168374 3060
rect 169450 2802 169478 3060
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 162814 2790 162866 2796
rect 163884 2774 163958 2802
rect 164988 2774 165062 2802
rect 166092 2774 166166 2802
rect 167196 2774 167270 2802
rect 168024 2774 168374 2802
rect 169404 2774 169478 2802
rect 156602 2408 156658 2417
rect 156602 2343 156658 2352
rect 156144 1352 156196 1358
rect 156144 1294 156196 1300
rect 156616 480 156644 2343
rect 158364 2009 158392 2774
rect 159468 2553 159496 2774
rect 160572 2689 160600 2774
rect 160558 2680 160614 2689
rect 160558 2615 160614 2624
rect 159454 2544 159510 2553
rect 159454 2479 159510 2488
rect 158350 2000 158406 2009
rect 158350 1935 158406 1944
rect 161294 2000 161350 2009
rect 161294 1935 161350 1944
rect 157798 1728 157854 1737
rect 157798 1663 157854 1672
rect 157812 480 157840 1663
rect 160112 598 160324 626
rect 160112 480 160140 598
rect 160296 513 160324 598
rect 160282 504 160338 513
rect 155040 196 155092 202
rect 155040 138 155092 144
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161308 480 161336 1935
rect 161676 1873 161704 2774
rect 162490 2544 162546 2553
rect 162490 2479 162546 2488
rect 161662 1864 161718 1873
rect 161662 1799 161718 1808
rect 162504 480 162532 2479
rect 163884 2145 163912 2774
rect 164988 2281 165016 2774
rect 166092 2417 166120 2774
rect 166078 2408 166134 2417
rect 166078 2343 166134 2352
rect 164974 2272 165030 2281
rect 164974 2207 165030 2216
rect 163870 2136 163926 2145
rect 163870 2071 163926 2080
rect 167196 1737 167224 2774
rect 167182 1728 167238 1737
rect 167182 1663 167238 1672
rect 164148 1352 164200 1358
rect 164148 1294 164200 1300
rect 164882 1320 164938 1329
rect 160282 439 160338 448
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 165908 377 165936 598
rect 166092 480 166120 598
rect 167196 480 167224 711
rect 165894 368 165950 377
rect 165894 303 165950 312
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169588 480 169616 2858
rect 170554 2802 170582 3060
rect 171658 2802 171686 3060
rect 172762 2802 172790 3060
rect 173866 2802 173894 3060
rect 174970 2802 174998 3060
rect 176074 2802 176102 3060
rect 177178 2802 177206 3060
rect 178282 2922 178310 3060
rect 178270 2916 178322 2922
rect 178270 2858 178322 2864
rect 179386 2802 179414 3060
rect 180490 2802 180518 3060
rect 181594 2802 181622 3060
rect 182698 2802 182726 3060
rect 183802 2802 183830 3060
rect 184906 2802 184934 3060
rect 186010 2802 186038 3060
rect 170508 2774 170582 2802
rect 171612 2774 171686 2802
rect 172716 2774 172790 2802
rect 173820 2774 173894 2802
rect 174924 2774 174998 2802
rect 176028 2774 176102 2802
rect 177132 2774 177206 2802
rect 179340 2774 179414 2802
rect 180444 2774 180518 2802
rect 181548 2774 181622 2802
rect 182652 2774 182726 2802
rect 183572 2774 183830 2802
rect 184860 2774 184934 2802
rect 185964 2774 186038 2802
rect 186134 2816 186190 2825
rect 170508 2009 170536 2774
rect 171612 2553 171640 2774
rect 171598 2544 171654 2553
rect 171598 2479 171654 2488
rect 170494 2000 170550 2009
rect 170494 1935 170550 1944
rect 172716 1358 172744 2774
rect 172704 1352 172756 1358
rect 173820 1329 173848 2774
rect 172704 1294 172756 1300
rect 173806 1320 173862 1329
rect 173806 1255 173862 1264
rect 174266 1320 174322 1329
rect 174266 1255 174322 1264
rect 171966 1184 172022 1193
rect 171966 1119 172022 1128
rect 170586 504 170642 513
rect 169390 439 169446 448
rect 169546 -960 169658 480
rect 171980 480 172008 1119
rect 173162 640 173218 649
rect 173162 575 173218 584
rect 173176 480 173204 575
rect 174280 480 174308 1255
rect 170586 439 170642 448
rect 170600 354 170628 439
rect 170742 354 170854 480
rect 170600 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 176856 377 176884 598
rect 177868 480 177896 983
rect 179050 776 179106 785
rect 179050 711 179106 720
rect 179064 480 179092 711
rect 179340 513 179368 2774
rect 180246 2000 180302 2009
rect 180246 1935 180302 1944
rect 179326 504 179382 513
rect 176842 368 176898 377
rect 176842 303 176898 312
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180260 480 180288 1935
rect 180444 1193 180472 2774
rect 180430 1184 180486 1193
rect 180430 1119 180486 1128
rect 181442 912 181498 921
rect 181442 847 181498 856
rect 181456 480 181484 847
rect 181548 649 181576 2774
rect 182652 1329 182680 2774
rect 182638 1320 182694 1329
rect 182638 1255 182694 1264
rect 181534 640 181590 649
rect 181534 575 181590 584
rect 179326 439 179382 448
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182362 232 182418 241
rect 182518 218 182630 480
rect 182418 190 182630 218
rect 182362 167 182418 176
rect 182518 -960 182630 190
rect 183466 96 183522 105
rect 183572 82 183600 2774
rect 183742 1184 183798 1193
rect 183742 1119 183798 1128
rect 183756 480 183784 1119
rect 184860 649 184888 2774
rect 184938 1320 184994 1329
rect 184938 1255 184994 1264
rect 184846 640 184902 649
rect 184846 575 184902 584
rect 184952 480 184980 1255
rect 185964 1057 185992 2774
rect 187114 2802 187142 3060
rect 188218 2802 188246 3060
rect 189322 2802 189350 3060
rect 190426 2802 190454 3060
rect 191530 2802 191558 3060
rect 192634 2802 192662 3060
rect 193738 2825 193766 3060
rect 186134 2751 186190 2760
rect 187068 2774 187142 2802
rect 188172 2774 188246 2802
rect 189276 2774 189350 2802
rect 190380 2774 190454 2802
rect 191484 2774 191558 2802
rect 192588 2774 192662 2802
rect 193724 2816 193780 2825
rect 185950 1048 186006 1057
rect 185950 983 186006 992
rect 186148 480 186176 2751
rect 187068 785 187096 2774
rect 188172 2009 188200 2774
rect 188158 2000 188214 2009
rect 188158 1935 188214 1944
rect 189276 921 189304 2774
rect 189722 2000 189778 2009
rect 189722 1935 189778 1944
rect 189262 912 189318 921
rect 189262 847 189318 856
rect 187054 776 187110 785
rect 187054 711 187110 720
rect 189736 480 189764 1935
rect 183522 54 183600 82
rect 183466 31 183522 40
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190380 241 190408 2774
rect 191484 1193 191512 2774
rect 192588 1329 192616 2774
rect 194842 2802 194870 3060
rect 195946 2802 195974 3060
rect 197050 2802 197078 3060
rect 198154 2802 198182 3060
rect 199258 2802 199286 3060
rect 200362 2802 200390 3060
rect 201466 2802 201494 3060
rect 202570 2802 202598 3060
rect 203674 2802 203702 3060
rect 204778 2802 204806 3060
rect 205882 2802 205910 3060
rect 206986 2802 207014 3060
rect 208090 2802 208118 3060
rect 209194 2802 209222 3060
rect 210298 2802 210326 3060
rect 211402 2802 211430 3060
rect 212506 2802 212534 3060
rect 213610 2802 213638 3060
rect 214714 2802 214742 3060
rect 215818 2802 215846 3060
rect 193724 2751 193780 2760
rect 194796 2774 194870 2802
rect 195900 2774 195974 2802
rect 197004 2774 197078 2802
rect 198108 2774 198182 2802
rect 199212 2774 199286 2802
rect 200316 2774 200390 2802
rect 201420 2774 201494 2802
rect 202524 2774 202598 2802
rect 203536 2774 203702 2802
rect 204732 2774 204806 2802
rect 205836 2774 205910 2802
rect 206940 2774 207014 2802
rect 208044 2774 208118 2802
rect 209148 2774 209222 2802
rect 210252 2774 210326 2802
rect 211356 2774 211430 2802
rect 212460 2774 212534 2802
rect 213564 2774 213638 2802
rect 214668 2774 214742 2802
rect 215772 2774 215846 2802
rect 216922 2802 216950 3060
rect 218026 2802 218054 3060
rect 219130 2802 219158 3060
rect 220234 2802 220262 3060
rect 221338 2802 221366 3060
rect 222442 2802 222470 3060
rect 223546 2802 223574 3060
rect 224650 2802 224678 3060
rect 225754 2802 225782 3060
rect 226858 2802 226886 3060
rect 227962 2802 227990 3060
rect 229066 2802 229094 3060
rect 230170 2802 230198 3060
rect 231274 2802 231302 3060
rect 232378 2802 232406 3060
rect 233482 2802 233510 3060
rect 234586 2802 234614 3060
rect 235690 2802 235718 3060
rect 236794 2802 236822 3060
rect 237898 2802 237926 3060
rect 239002 2802 239030 3060
rect 240106 2802 240134 3060
rect 241210 2802 241238 3060
rect 242314 2802 242342 3060
rect 243418 2802 243446 3060
rect 244522 2802 244550 3060
rect 245626 2802 245654 3060
rect 246730 2802 246758 3060
rect 247834 2802 247862 3060
rect 248938 2802 248966 3060
rect 250042 2802 250070 3060
rect 251146 2802 251174 3060
rect 252250 2802 252278 3060
rect 253354 2802 253382 3060
rect 254458 2802 254486 3060
rect 255562 2802 255590 3060
rect 256666 2802 256694 3060
rect 257770 2802 257798 3060
rect 258874 2802 258902 3060
rect 259978 2802 260006 3060
rect 261082 2802 261110 3060
rect 262186 2802 262214 3060
rect 263290 2802 263318 3060
rect 264394 2802 264422 3060
rect 265498 2802 265526 3060
rect 266602 2802 266630 3060
rect 267706 2802 267734 3060
rect 268810 2802 268838 3060
rect 269914 2802 269942 3060
rect 271018 2802 271046 3060
rect 272122 2802 272150 3060
rect 273226 2802 273254 3060
rect 274330 2802 274358 3060
rect 275434 2802 275462 3060
rect 276538 2802 276566 3060
rect 277642 2802 277670 3060
rect 278746 2802 278774 3060
rect 279850 2802 279878 3060
rect 280954 2802 280982 3060
rect 282058 2802 282086 3060
rect 283162 2938 283190 3060
rect 284266 2938 284294 3060
rect 283162 2910 283236 2938
rect 216922 2774 216996 2802
rect 192574 1320 192630 1329
rect 192574 1255 192630 1264
rect 191470 1184 191526 1193
rect 191470 1119 191526 1128
rect 194414 1184 194470 1193
rect 194414 1119 194470 1128
rect 193218 1048 193274 1057
rect 193218 983 193274 992
rect 192022 912 192078 921
rect 192022 847 192078 856
rect 190826 776 190882 785
rect 190826 711 190882 720
rect 190840 480 190868 711
rect 192036 480 192064 847
rect 193232 480 193260 983
rect 194428 480 194456 1119
rect 190366 232 190422 241
rect 190366 167 190422 176
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 194796 105 194824 2774
rect 195610 1320 195666 1329
rect 195610 1255 195666 1264
rect 195624 480 195652 1255
rect 195900 649 195928 2774
rect 197004 2009 197032 2774
rect 196990 2000 197046 2009
rect 196990 1935 197046 1944
rect 198108 785 198136 2774
rect 199212 921 199240 2774
rect 200316 1057 200344 2774
rect 200486 1728 200542 1737
rect 200408 1686 200486 1714
rect 200302 1048 200358 1057
rect 200302 983 200358 992
rect 199198 912 199254 921
rect 200408 898 200436 1686
rect 200486 1663 200542 1672
rect 201420 1193 201448 2774
rect 201498 1456 201554 1465
rect 201498 1391 201554 1400
rect 201406 1184 201462 1193
rect 201406 1119 201462 1128
rect 199198 847 199254 856
rect 200316 870 200436 898
rect 198094 776 198150 785
rect 198094 711 198150 720
rect 199106 776 199162 785
rect 199106 711 199162 720
rect 195886 640 195942 649
rect 195886 575 195942 584
rect 199120 480 199148 711
rect 200316 480 200344 870
rect 201512 480 201540 1391
rect 202524 1329 202552 2774
rect 202510 1320 202566 1329
rect 202510 1255 202566 1264
rect 202694 1048 202750 1057
rect 202694 983 202750 992
rect 202708 480 202736 983
rect 194782 96 194838 105
rect 194782 31 194838 40
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203536 105 203564 2774
rect 203890 1184 203946 1193
rect 203890 1119 203946 1128
rect 203904 480 203932 1119
rect 203522 96 203578 105
rect 203522 31 203578 40
rect 203862 -960 203974 480
rect 204732 377 204760 2774
rect 205086 1320 205142 1329
rect 205086 1255 205142 1264
rect 205100 480 205128 1255
rect 205836 785 205864 2774
rect 206940 1737 206968 2774
rect 207386 2136 207442 2145
rect 207386 2071 207442 2080
rect 206926 1728 206982 1737
rect 206926 1663 206982 1672
rect 206190 1592 206246 1601
rect 206190 1527 206246 1536
rect 205822 776 205878 785
rect 205822 711 205878 720
rect 206204 480 206232 1527
rect 207400 480 207428 2071
rect 208044 1465 208072 2774
rect 208582 2000 208638 2009
rect 208582 1935 208638 1944
rect 208030 1456 208086 1465
rect 208030 1391 208086 1400
rect 208596 480 208624 1935
rect 209148 1057 209176 2774
rect 209778 2272 209834 2281
rect 209778 2207 209834 2216
rect 209134 1048 209190 1057
rect 209134 983 209190 992
rect 209792 480 209820 2207
rect 210252 1193 210280 2774
rect 211356 1329 211384 2774
rect 212170 1864 212226 1873
rect 212170 1799 212226 1808
rect 211342 1320 211398 1329
rect 211342 1255 211398 1264
rect 210238 1184 210294 1193
rect 210238 1119 210294 1128
rect 210974 1184 211030 1193
rect 210974 1119 211030 1128
rect 210988 480 211016 1119
rect 212184 480 212212 1799
rect 212460 1601 212488 2774
rect 213564 2145 213592 2774
rect 213550 2136 213606 2145
rect 213550 2071 213606 2080
rect 214668 2009 214696 2774
rect 215772 2281 215800 2774
rect 216862 2408 216918 2417
rect 216862 2343 216918 2352
rect 215758 2272 215814 2281
rect 215758 2207 215814 2216
rect 214654 2000 214710 2009
rect 214654 1935 214710 1944
rect 213366 1728 213422 1737
rect 213366 1663 213422 1672
rect 212446 1592 212502 1601
rect 212446 1527 212502 1536
rect 213380 480 213408 1663
rect 215666 1592 215722 1601
rect 215666 1527 215722 1536
rect 214470 1456 214526 1465
rect 214470 1391 214526 1400
rect 214484 480 214512 1391
rect 215680 480 215708 1527
rect 216876 480 216904 2343
rect 216968 1193 216996 2774
rect 217980 2774 218054 2802
rect 219084 2774 219158 2802
rect 220188 2774 220262 2802
rect 221292 2774 221366 2802
rect 222396 2774 222470 2802
rect 223500 2774 223574 2802
rect 224604 2774 224678 2802
rect 225708 2774 225782 2802
rect 226812 2774 226886 2802
rect 227916 2774 227990 2802
rect 229020 2774 229094 2802
rect 230124 2774 230198 2802
rect 231228 2774 231302 2802
rect 232332 2774 232406 2802
rect 233436 2774 233510 2802
rect 234540 2774 234614 2802
rect 235644 2774 235718 2802
rect 236748 2774 236822 2802
rect 237852 2774 237926 2802
rect 238956 2774 239030 2802
rect 240060 2774 240134 2802
rect 241164 2774 241238 2802
rect 242268 2774 242342 2802
rect 243372 2774 243446 2802
rect 244476 2774 244550 2802
rect 245580 2774 245654 2802
rect 246684 2774 246758 2802
rect 247788 2774 247862 2802
rect 248892 2774 248966 2802
rect 249996 2774 250070 2802
rect 251100 2774 251174 2802
rect 252204 2774 252278 2802
rect 253308 2774 253382 2802
rect 254412 2774 254486 2802
rect 255516 2774 255590 2802
rect 256620 2774 256694 2802
rect 257724 2774 257798 2802
rect 258828 2774 258902 2802
rect 259932 2774 260006 2802
rect 261036 2774 261110 2802
rect 262140 2774 262214 2802
rect 263244 2774 263318 2802
rect 264348 2774 264422 2802
rect 265452 2774 265526 2802
rect 266556 2774 266630 2802
rect 267660 2774 267734 2802
rect 268764 2774 268838 2802
rect 269868 2774 269942 2802
rect 270972 2774 271046 2802
rect 272076 2774 272150 2802
rect 273180 2774 273254 2802
rect 274284 2774 274358 2802
rect 275388 2774 275462 2802
rect 276492 2774 276566 2802
rect 277596 2774 277670 2802
rect 278700 2774 278774 2802
rect 279804 2774 279878 2802
rect 280908 2774 280982 2802
rect 282012 2774 282086 2802
rect 217980 1873 218008 2774
rect 218058 2680 218114 2689
rect 218058 2615 218114 2624
rect 217966 1864 218022 1873
rect 217966 1799 218022 1808
rect 216954 1184 217010 1193
rect 216954 1119 217010 1128
rect 218072 480 218100 2615
rect 219084 1737 219112 2774
rect 219254 2272 219310 2281
rect 219254 2207 219310 2216
rect 219070 1728 219126 1737
rect 219070 1663 219126 1672
rect 219268 480 219296 2207
rect 220188 1465 220216 2774
rect 220450 2000 220506 2009
rect 220450 1935 220506 1944
rect 220174 1456 220230 1465
rect 220174 1391 220230 1400
rect 220464 480 220492 1935
rect 221292 1601 221320 2774
rect 222396 2417 222424 2774
rect 223500 2689 223528 2774
rect 223486 2680 223542 2689
rect 223486 2615 223542 2624
rect 222382 2408 222438 2417
rect 222382 2343 222438 2352
rect 224604 2281 224632 2774
rect 224590 2272 224646 2281
rect 224590 2207 224646 2216
rect 223946 2136 224002 2145
rect 223946 2071 224002 2080
rect 221554 1864 221610 1873
rect 221554 1799 221610 1808
rect 221278 1592 221334 1601
rect 221278 1527 221334 1536
rect 221568 480 221596 1799
rect 222750 1728 222806 1737
rect 222750 1663 222806 1672
rect 222764 480 222792 1663
rect 223960 480 223988 2071
rect 225708 2009 225736 2774
rect 225694 2000 225750 2009
rect 225694 1935 225750 1944
rect 226812 1873 226840 2774
rect 227534 2000 227590 2009
rect 227534 1935 227590 1944
rect 226798 1864 226854 1873
rect 226798 1799 226854 1808
rect 226338 1592 226394 1601
rect 226338 1527 226394 1536
rect 225142 1456 225198 1465
rect 225142 1391 225198 1400
rect 225156 480 225184 1391
rect 226352 480 226380 1527
rect 227548 480 227576 1935
rect 227916 1737 227944 2774
rect 228730 2408 228786 2417
rect 228730 2343 228786 2352
rect 227902 1728 227958 1737
rect 227902 1663 227958 1672
rect 228744 480 228772 2343
rect 229020 2145 229048 2774
rect 229006 2136 229062 2145
rect 229006 2071 229062 2080
rect 229834 2136 229890 2145
rect 229834 2071 229890 2080
rect 229848 480 229876 2071
rect 230124 1465 230152 2774
rect 231228 1601 231256 2774
rect 232332 2009 232360 2774
rect 233436 2417 233464 2774
rect 233422 2408 233478 2417
rect 233422 2343 233478 2352
rect 234540 2145 234568 2774
rect 234526 2136 234582 2145
rect 234526 2071 234582 2080
rect 232318 2000 232374 2009
rect 232318 1935 232374 1944
rect 233422 1864 233478 1873
rect 233422 1799 233478 1808
rect 231214 1592 231270 1601
rect 231214 1527 231270 1536
rect 232226 1592 232282 1601
rect 232226 1527 232282 1536
rect 230110 1456 230166 1465
rect 230110 1391 230166 1400
rect 231030 1456 231086 1465
rect 231030 1391 231086 1400
rect 231044 480 231072 1391
rect 232240 480 232268 1527
rect 233436 480 233464 1799
rect 234618 1728 234674 1737
rect 234618 1663 234674 1672
rect 234632 480 234660 1663
rect 235644 1465 235672 2774
rect 236748 1601 236776 2774
rect 237852 1873 237880 2774
rect 238114 2000 238170 2009
rect 238114 1935 238170 1944
rect 237838 1864 237894 1873
rect 237838 1799 237894 1808
rect 236734 1592 236790 1601
rect 236734 1527 236790 1536
rect 237010 1592 237066 1601
rect 237010 1527 237066 1536
rect 235630 1456 235686 1465
rect 235630 1391 235686 1400
rect 235814 1456 235870 1465
rect 235814 1391 235870 1400
rect 235828 480 235856 1391
rect 237024 480 237052 1527
rect 238128 480 238156 1935
rect 238956 1737 238984 2774
rect 239310 2136 239366 2145
rect 239310 2071 239366 2080
rect 238942 1728 238998 1737
rect 238942 1663 238998 1672
rect 239324 480 239352 2071
rect 240060 1465 240088 2774
rect 241164 1601 241192 2774
rect 242268 2009 242296 2774
rect 243372 2145 243400 2774
rect 243358 2136 243414 2145
rect 243358 2071 243414 2080
rect 242254 2000 242310 2009
rect 242254 1935 242310 1944
rect 241702 1864 241758 1873
rect 241702 1799 241758 1808
rect 241150 1592 241206 1601
rect 241150 1527 241206 1536
rect 240046 1456 240102 1465
rect 240046 1391 240102 1400
rect 240506 1456 240562 1465
rect 240506 1391 240562 1400
rect 240520 480 240548 1391
rect 241716 480 241744 1799
rect 242898 1728 242954 1737
rect 242898 1663 242954 1672
rect 242912 480 242940 1663
rect 244094 1592 244150 1601
rect 244094 1527 244150 1536
rect 244108 480 244136 1527
rect 244476 1465 244504 2774
rect 245580 1873 245608 2774
rect 246394 2408 246450 2417
rect 246394 2343 246450 2352
rect 245566 1864 245622 1873
rect 245566 1799 245622 1808
rect 244462 1456 244518 1465
rect 244462 1391 244518 1400
rect 245198 1456 245254 1465
rect 245198 1391 245254 1400
rect 245212 480 245240 1391
rect 246408 480 246436 2343
rect 246684 1737 246712 2774
rect 247590 1864 247646 1873
rect 247590 1799 247646 1808
rect 246670 1728 246726 1737
rect 246670 1663 246726 1672
rect 247604 480 247632 1799
rect 247788 1601 247816 2774
rect 248786 2000 248842 2009
rect 248786 1935 248842 1944
rect 247774 1592 247830 1601
rect 247774 1527 247830 1536
rect 248800 480 248828 1935
rect 248892 1465 248920 2774
rect 249996 2417 250024 2774
rect 249982 2408 250038 2417
rect 249982 2343 250038 2352
rect 251100 1873 251128 2774
rect 252204 2009 252232 2774
rect 252190 2000 252246 2009
rect 252190 1935 252246 1944
rect 251086 1864 251142 1873
rect 251086 1799 251142 1808
rect 251178 1728 251234 1737
rect 251178 1663 251234 1672
rect 249982 1592 250038 1601
rect 249982 1527 250038 1536
rect 248878 1456 248934 1465
rect 248878 1391 248934 1400
rect 249996 480 250024 1527
rect 251192 480 251220 1663
rect 253308 1601 253336 2774
rect 254412 1737 254440 2774
rect 254398 1728 254454 1737
rect 254398 1663 254454 1672
rect 254674 1728 254730 1737
rect 254674 1663 254730 1672
rect 253294 1592 253350 1601
rect 253294 1527 253350 1536
rect 253478 1592 253534 1601
rect 253478 1527 253534 1536
rect 252374 1456 252430 1465
rect 252374 1391 252430 1400
rect 252388 480 252416 1391
rect 253492 480 253520 1527
rect 254688 480 254716 1663
rect 255516 1465 255544 2774
rect 256620 1601 256648 2774
rect 257724 1737 257752 2774
rect 257710 1728 257766 1737
rect 257710 1663 257766 1672
rect 258262 1728 258318 1737
rect 258262 1663 258318 1672
rect 256606 1592 256662 1601
rect 256606 1527 256662 1536
rect 257066 1592 257122 1601
rect 257066 1527 257122 1536
rect 255502 1456 255558 1465
rect 255502 1391 255558 1400
rect 255870 1456 255926 1465
rect 255870 1391 255926 1400
rect 255884 480 255912 1391
rect 257080 480 257108 1527
rect 258276 480 258304 1663
rect 258828 1465 258856 2774
rect 259932 1601 259960 2774
rect 261036 1737 261064 2774
rect 261022 1728 261078 1737
rect 261022 1663 261078 1672
rect 261758 1728 261814 1737
rect 261758 1663 261814 1672
rect 259918 1592 259974 1601
rect 259918 1527 259974 1536
rect 260654 1592 260710 1601
rect 260654 1527 260710 1536
rect 258814 1456 258870 1465
rect 258814 1391 258870 1400
rect 259458 1320 259514 1329
rect 259458 1255 259514 1264
rect 259472 480 259500 1255
rect 260668 480 260696 1527
rect 261772 480 261800 1663
rect 262140 1329 262168 2774
rect 263244 1601 263272 2774
rect 264348 1737 264376 2774
rect 264334 1728 264390 1737
rect 264334 1663 264390 1672
rect 263230 1592 263286 1601
rect 263230 1527 263286 1536
rect 264150 1592 264206 1601
rect 264150 1527 264206 1536
rect 262954 1456 263010 1465
rect 262954 1391 263010 1400
rect 262126 1320 262182 1329
rect 262126 1255 262182 1264
rect 262968 480 262996 1391
rect 264164 480 264192 1527
rect 265452 1465 265480 2774
rect 266556 1601 266584 2774
rect 266542 1592 266598 1601
rect 266542 1527 266598 1536
rect 265438 1456 265494 1465
rect 265438 1391 265494 1400
rect 266542 1184 266598 1193
rect 266542 1119 266598 1128
rect 265346 1048 265402 1057
rect 265346 983 265402 992
rect 265360 480 265388 983
rect 266556 480 266584 1119
rect 267660 1057 267688 2774
rect 267738 1320 267794 1329
rect 267738 1255 267794 1264
rect 267646 1048 267702 1057
rect 267646 983 267702 992
rect 267752 480 267780 1255
rect 268764 1193 268792 2774
rect 268842 1456 268898 1465
rect 268842 1391 268898 1400
rect 268750 1184 268806 1193
rect 268750 1119 268806 1128
rect 268856 480 268884 1391
rect 269868 1329 269896 2774
rect 270038 1592 270094 1601
rect 270038 1527 270094 1536
rect 269854 1320 269910 1329
rect 269854 1255 269910 1264
rect 270052 480 270080 1527
rect 270972 1465 271000 2774
rect 272076 1601 272104 2774
rect 272062 1592 272118 1601
rect 272062 1527 272118 1536
rect 270958 1456 271014 1465
rect 270958 1391 271014 1400
rect 273180 1329 273208 2774
rect 271234 1320 271290 1329
rect 271234 1255 271290 1264
rect 273166 1320 273222 1329
rect 273166 1255 273222 1264
rect 273626 1320 273682 1329
rect 273626 1255 273682 1264
rect 271248 480 271276 1255
rect 272430 1184 272486 1193
rect 272430 1119 272486 1128
rect 272444 480 272472 1119
rect 273640 480 273668 1255
rect 274284 1193 274312 2774
rect 275388 1329 275416 2774
rect 275374 1320 275430 1329
rect 275374 1255 275430 1264
rect 276018 1320 276074 1329
rect 276018 1255 276074 1264
rect 274270 1184 274326 1193
rect 274270 1119 274326 1128
rect 274822 1184 274878 1193
rect 274822 1119 274878 1128
rect 274836 480 274864 1119
rect 276032 480 276060 1255
rect 276492 1193 276520 2774
rect 277596 1329 277624 2774
rect 277582 1320 277638 1329
rect 277582 1255 277638 1264
rect 278700 1193 278728 2774
rect 279514 1320 279570 1329
rect 279514 1255 279570 1264
rect 276478 1184 276534 1193
rect 276478 1119 276534 1128
rect 277122 1184 277178 1193
rect 277122 1119 277178 1128
rect 278686 1184 278742 1193
rect 278686 1119 278742 1128
rect 277136 480 277164 1119
rect 278318 1048 278374 1057
rect 278318 983 278374 992
rect 278332 480 278360 983
rect 279528 480 279556 1255
rect 279804 1057 279832 2774
rect 280908 1329 280936 2774
rect 280894 1320 280950 1329
rect 280894 1255 280950 1264
rect 281906 1320 281962 1329
rect 281906 1255 281962 1264
rect 280710 1184 280766 1193
rect 280710 1119 280766 1128
rect 279790 1048 279846 1057
rect 279790 983 279846 992
rect 280724 480 280752 1119
rect 281920 480 281948 1255
rect 282012 1193 282040 2774
rect 283208 1329 283236 2910
rect 283300 2910 284294 2938
rect 283194 1320 283250 1329
rect 283194 1255 283250 1264
rect 281998 1184 282054 1193
rect 283300 1170 283328 2910
rect 285370 2802 285398 3060
rect 286474 2802 286502 3060
rect 287578 2802 287606 3060
rect 288682 2802 288710 3060
rect 289786 2802 289814 3060
rect 290890 2802 290918 3060
rect 291994 2802 292022 3060
rect 293098 2802 293126 3060
rect 294202 2802 294230 3060
rect 295306 2802 295334 3060
rect 296410 2802 296438 3060
rect 297514 2802 297542 3060
rect 298618 2802 298646 3060
rect 299722 2802 299750 3060
rect 300826 2802 300854 3060
rect 281998 1119 282054 1128
rect 283116 1142 283328 1170
rect 284312 2774 285398 2802
rect 286428 2774 286502 2802
rect 287532 2774 287606 2802
rect 288636 2774 288710 2802
rect 289464 2774 289814 2802
rect 290200 2774 290918 2802
rect 291856 2774 292022 2802
rect 292592 2774 293126 2802
rect 293696 2774 294230 2802
rect 295260 2774 295334 2802
rect 296088 2774 296438 2802
rect 297468 2774 297542 2802
rect 298480 2774 298646 2802
rect 299676 2774 299750 2802
rect 300780 2774 300854 2802
rect 301930 2802 301958 3060
rect 303034 2802 303062 3060
rect 304138 2802 304166 3060
rect 305242 2802 305270 3060
rect 306346 2802 306374 3060
rect 307450 2802 307478 3060
rect 308554 2802 308582 3060
rect 309658 2802 309686 3060
rect 310762 2802 310790 3060
rect 311866 2802 311894 3060
rect 312970 2802 312998 3060
rect 314074 2802 314102 3060
rect 315178 2802 315206 3060
rect 316282 2802 316310 3060
rect 317386 2938 317414 3060
rect 317386 2910 317460 2938
rect 301930 2774 302004 2802
rect 303034 2774 303200 2802
rect 304138 2774 304212 2802
rect 305242 2774 305592 2802
rect 306346 2774 306420 2802
rect 307450 2774 307984 2802
rect 308554 2774 309088 2802
rect 309658 2774 309824 2802
rect 310762 2774 311480 2802
rect 311866 2774 312216 2802
rect 312970 2774 313044 2802
rect 314074 2774 314148 2802
rect 315178 2774 315252 2802
rect 316282 2774 317368 2802
rect 283116 480 283144 1142
rect 284312 480 284340 2774
rect 286428 1329 286456 2774
rect 287532 1329 287560 2774
rect 288636 1329 288664 2774
rect 285402 1320 285458 1329
rect 285402 1255 285458 1264
rect 286414 1320 286470 1329
rect 286414 1255 286470 1264
rect 286598 1320 286654 1329
rect 286598 1255 286654 1264
rect 287518 1320 287574 1329
rect 287518 1255 287574 1264
rect 287794 1320 287850 1329
rect 287794 1255 287850 1264
rect 288622 1320 288678 1329
rect 288622 1255 288678 1264
rect 285416 480 285444 1255
rect 286612 480 286640 1255
rect 287808 480 287836 1255
rect 204718 368 204774 377
rect 204718 303 204774 312
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289464 354 289492 2774
rect 290200 480 290228 2774
rect 288962 326 289492 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 354 291466 480
rect 291856 354 291884 2774
rect 292592 480 292620 2774
rect 293696 480 293724 2774
rect 291354 326 291884 354
rect 291354 -960 291466 326
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 354 294962 480
rect 295260 354 295288 2774
rect 296088 480 296116 2774
rect 294850 326 295288 354
rect 294850 -960 294962 326
rect 296046 -960 296158 480
rect 297242 354 297354 480
rect 297468 354 297496 2774
rect 298480 480 298508 2774
rect 299676 480 299704 2774
rect 300780 480 300808 2774
rect 301976 480 302004 2774
rect 303172 480 303200 2774
rect 297242 326 297496 354
rect 297242 -960 297354 326
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304184 354 304212 2774
rect 305564 480 305592 2774
rect 304326 354 304438 480
rect 304184 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 2774
rect 307956 480 307984 2774
rect 309060 480 309088 2774
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 2774
rect 311452 480 311480 2774
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 2774
rect 313016 1329 313044 2774
rect 314120 1329 314148 2774
rect 315224 1329 315252 2774
rect 313002 1320 313058 1329
rect 313002 1255 313058 1264
rect 313830 1320 313886 1329
rect 313830 1255 313886 1264
rect 314106 1320 314162 1329
rect 314106 1255 314162 1264
rect 315026 1320 315082 1329
rect 315026 1255 315082 1264
rect 315210 1320 315266 1329
rect 315210 1255 315266 1264
rect 316222 1320 316278 1329
rect 316222 1255 316278 1264
rect 313844 480 313872 1255
rect 315040 480 315068 1255
rect 316236 480 316264 1255
rect 317340 480 317368 2774
rect 317432 1329 317460 2910
rect 318490 2802 318518 3060
rect 318444 2774 318518 2802
rect 319594 2802 319622 3060
rect 320698 2802 320726 3060
rect 321802 2802 321830 3060
rect 322906 2802 322934 3060
rect 319594 2774 319668 2802
rect 320698 2774 320772 2802
rect 321802 2774 321876 2802
rect 317418 1320 317474 1329
rect 317418 1255 317474 1264
rect 318444 1193 318472 2774
rect 319640 1329 319668 2774
rect 318522 1320 318578 1329
rect 318522 1255 318578 1264
rect 319626 1320 319682 1329
rect 319626 1255 319682 1264
rect 318430 1184 318486 1193
rect 318430 1119 318486 1128
rect 318536 480 318564 1255
rect 320744 1193 320772 2774
rect 320914 1320 320970 1329
rect 320914 1255 320970 1264
rect 319718 1184 319774 1193
rect 319718 1119 319774 1128
rect 320730 1184 320786 1193
rect 320730 1119 320786 1128
rect 319732 480 319760 1119
rect 320928 480 320956 1255
rect 321848 1057 321876 2774
rect 322860 2774 322934 2802
rect 324010 2802 324038 3060
rect 325114 2802 325142 3060
rect 326218 2802 326246 3060
rect 327322 2802 327350 3060
rect 328426 2802 328454 3060
rect 324010 2774 324084 2802
rect 325114 2774 325188 2802
rect 326218 2774 326292 2802
rect 327322 2774 327396 2802
rect 322860 1329 322888 2774
rect 322846 1320 322902 1329
rect 322846 1255 322902 1264
rect 324056 1193 324084 2774
rect 325160 1329 325188 2774
rect 324410 1320 324466 1329
rect 324410 1255 324466 1264
rect 325146 1320 325202 1329
rect 325146 1255 325202 1264
rect 322110 1184 322166 1193
rect 322110 1119 322166 1128
rect 324042 1184 324098 1193
rect 324042 1119 324098 1128
rect 321834 1048 321890 1057
rect 321834 983 321890 992
rect 322124 480 322152 1119
rect 323306 1048 323362 1057
rect 323306 983 323362 992
rect 323320 480 323348 983
rect 324424 480 324452 1255
rect 326264 1193 326292 2774
rect 327368 1329 327396 2774
rect 328380 2774 328454 2802
rect 329530 2802 329558 3060
rect 330634 2802 330662 3060
rect 331738 2802 331766 3060
rect 332842 2802 332870 3060
rect 333946 2802 333974 3060
rect 329530 2774 329604 2802
rect 330634 2774 330708 2802
rect 331738 2774 331812 2802
rect 332842 2774 332916 2802
rect 326802 1320 326858 1329
rect 326802 1255 326858 1264
rect 327354 1320 327410 1329
rect 327354 1255 327410 1264
rect 325606 1184 325662 1193
rect 325606 1119 325662 1128
rect 326250 1184 326306 1193
rect 326250 1119 326306 1128
rect 325620 480 325648 1119
rect 326816 480 326844 1255
rect 328380 1193 328408 2774
rect 329576 1329 329604 2774
rect 329194 1320 329250 1329
rect 329194 1255 329250 1264
rect 329562 1320 329618 1329
rect 329562 1255 329618 1264
rect 327998 1184 328054 1193
rect 327998 1119 328054 1128
rect 328366 1184 328422 1193
rect 328366 1119 328422 1128
rect 328012 480 328040 1119
rect 329208 480 329236 1255
rect 330680 1193 330708 2774
rect 331586 1320 331642 1329
rect 331586 1255 331642 1264
rect 330390 1184 330446 1193
rect 330390 1119 330446 1128
rect 330666 1184 330722 1193
rect 330666 1119 330722 1128
rect 330404 480 330432 1119
rect 331600 480 331628 1255
rect 331784 921 331812 2774
rect 332888 1193 332916 2774
rect 333900 2774 333974 2802
rect 335050 2802 335078 3060
rect 336154 2802 336182 3060
rect 337258 2802 337286 3060
rect 338362 2802 338390 3060
rect 339466 2802 339494 3060
rect 335050 2774 335124 2802
rect 336154 2774 336228 2802
rect 337258 2774 337332 2802
rect 338362 2774 338436 2802
rect 332690 1184 332746 1193
rect 332690 1119 332746 1128
rect 332874 1184 332930 1193
rect 332874 1119 332930 1128
rect 331770 912 331826 921
rect 331770 847 331826 856
rect 332704 480 332732 1119
rect 333900 1057 333928 2774
rect 335096 1329 335124 2774
rect 335082 1320 335138 1329
rect 335082 1255 335138 1264
rect 336200 1193 336228 2774
rect 335082 1184 335138 1193
rect 335082 1119 335138 1128
rect 336186 1184 336242 1193
rect 336186 1119 336242 1128
rect 333886 1048 333942 1057
rect 333886 983 333942 992
rect 333886 912 333942 921
rect 333886 847 333942 856
rect 333900 480 333928 847
rect 335096 480 335124 1119
rect 337304 1057 337332 2774
rect 338408 1329 338436 2774
rect 339420 2774 339494 2802
rect 340570 2802 340598 3060
rect 341674 2802 341702 3060
rect 342778 2802 342806 3060
rect 343882 2802 343910 3060
rect 344986 2825 345014 3060
rect 346090 2825 346118 3060
rect 344972 2816 345028 2825
rect 340570 2774 340644 2802
rect 341674 2774 341748 2802
rect 342778 2774 342852 2802
rect 343882 2774 343956 2802
rect 337474 1320 337530 1329
rect 337474 1255 337530 1264
rect 338394 1320 338450 1329
rect 338394 1255 338450 1264
rect 336278 1048 336334 1057
rect 336278 983 336334 992
rect 337290 1048 337346 1057
rect 337290 983 337346 992
rect 336292 480 336320 983
rect 337488 480 337516 1255
rect 339420 1193 339448 2774
rect 338670 1184 338726 1193
rect 338670 1119 338726 1128
rect 339406 1184 339462 1193
rect 339406 1119 339462 1128
rect 338684 480 338712 1119
rect 340616 1057 340644 2774
rect 341720 1329 341748 2774
rect 340970 1320 341026 1329
rect 340970 1255 341026 1264
rect 341706 1320 341762 1329
rect 341706 1255 341762 1264
rect 339866 1048 339922 1057
rect 339866 983 339922 992
rect 340602 1048 340658 1057
rect 340602 983 340658 992
rect 339880 480 339908 983
rect 340984 480 341012 1255
rect 342824 1193 342852 2774
rect 342166 1184 342222 1193
rect 342166 1119 342222 1128
rect 342810 1184 342866 1193
rect 342810 1119 342866 1128
rect 342180 480 342208 1119
rect 343928 1057 343956 2774
rect 344972 2751 345028 2760
rect 346076 2816 346132 2825
rect 347194 2802 347222 3060
rect 348298 2802 348326 3060
rect 349250 2816 349306 2825
rect 347194 2774 347268 2802
rect 348298 2774 348372 2802
rect 346076 2751 346132 2760
rect 347240 1329 347268 2774
rect 347778 2680 347834 2689
rect 347834 2638 348096 2666
rect 347778 2615 347834 2624
rect 344558 1320 344614 1329
rect 344558 1255 344614 1264
rect 347226 1320 347282 1329
rect 347226 1255 347282 1264
rect 343362 1048 343418 1057
rect 343362 983 343418 992
rect 343914 1048 343970 1057
rect 343914 983 343970 992
rect 343376 480 343404 983
rect 344572 480 344600 1255
rect 345754 1184 345810 1193
rect 345754 1119 345810 1128
rect 345768 480 345796 1119
rect 346950 1048 347006 1057
rect 346950 983 347006 992
rect 346964 480 346992 983
rect 348068 480 348096 2638
rect 348344 1193 348372 2774
rect 349402 2802 349430 3060
rect 350506 2825 350534 3060
rect 351610 2854 351638 3060
rect 351598 2848 351650 2854
rect 350492 2816 350548 2825
rect 349402 2774 349476 2802
rect 349250 2751 349306 2760
rect 348330 1184 348386 1193
rect 348330 1119 348386 1128
rect 349264 480 349292 2751
rect 349448 1057 349476 2774
rect 352714 2825 352742 3060
rect 353818 2961 353846 3060
rect 353804 2952 353860 2961
rect 353804 2887 353860 2896
rect 351598 2790 351650 2796
rect 352700 2816 352756 2825
rect 350492 2751 350548 2760
rect 354922 2802 354950 3060
rect 355048 2848 355100 2854
rect 354922 2774 354996 2802
rect 355048 2790 355100 2796
rect 356026 2802 356054 3060
rect 357130 2825 357158 3060
rect 358234 2854 358262 3060
rect 359338 2922 359366 3060
rect 360442 2961 360470 3060
rect 360428 2952 360484 2961
rect 359326 2916 359378 2922
rect 360428 2887 360484 2896
rect 359326 2858 359378 2864
rect 358222 2848 358274 2854
rect 356334 2816 356390 2825
rect 352700 2751 352756 2760
rect 353298 2680 353354 2689
rect 353354 2638 353616 2666
rect 353298 2615 353354 2624
rect 350446 1320 350502 1329
rect 350446 1255 350502 1264
rect 349434 1048 349490 1057
rect 349434 983 349490 992
rect 350460 480 350488 1255
rect 351642 1184 351698 1193
rect 351642 1119 351698 1128
rect 351656 480 351684 1119
rect 352838 1048 352894 1057
rect 352838 983 352894 992
rect 352852 480 352880 983
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 2638
rect 354968 1329 354996 2774
rect 355060 1442 355088 2790
rect 356026 2774 356100 2802
rect 356072 2689 356100 2774
rect 356334 2751 356390 2760
rect 356886 2816 356942 2825
rect 357116 2816 357172 2825
rect 356942 2774 357020 2802
rect 356886 2751 356942 2760
rect 356058 2680 356114 2689
rect 356058 2615 356114 2624
rect 355060 1414 355272 1442
rect 354954 1320 355010 1329
rect 354954 1255 355010 1264
rect 355244 480 355272 1414
rect 356348 480 356376 2751
rect 356992 2666 357020 2774
rect 361546 2825 361574 3060
rect 361672 2848 361724 2854
rect 358222 2790 358274 2796
rect 359922 2816 359978 2825
rect 357116 2751 357172 2760
rect 359922 2751 359978 2760
rect 361118 2816 361174 2825
rect 361118 2751 361174 2760
rect 361532 2816 361588 2825
rect 362650 2802 362678 3060
rect 363754 2961 363782 3060
rect 363740 2952 363796 2961
rect 363328 2916 363380 2922
rect 363740 2887 363796 2896
rect 364064 2916 364116 2922
rect 363328 2858 363380 2864
rect 364064 2858 364116 2864
rect 361724 2796 361896 2802
rect 361672 2790 361896 2796
rect 361684 2774 361896 2790
rect 362650 2774 362724 2802
rect 361532 2751 361588 2760
rect 356992 2638 357572 2666
rect 357544 480 357572 2638
rect 358726 1320 358782 1329
rect 358726 1255 358782 1264
rect 358740 480 358768 1255
rect 359936 480 359964 2751
rect 361132 480 361160 2751
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 2774
rect 362696 1562 362724 2774
rect 363340 1578 363368 2858
rect 364076 2825 364104 2858
rect 364858 2825 364886 3060
rect 365962 2922 365990 3060
rect 365720 2916 365772 2922
rect 365720 2858 365772 2864
rect 365950 2916 366002 2922
rect 365950 2858 366002 2864
rect 364062 2816 364118 2825
rect 364062 2751 364118 2760
rect 364614 2816 364670 2825
rect 364614 2751 364670 2760
rect 364844 2816 364900 2825
rect 364844 2751 364900 2760
rect 362684 1556 362736 1562
rect 363340 1550 363552 1578
rect 362684 1498 362736 1504
rect 363524 480 363552 1550
rect 364628 480 364656 2751
rect 365732 1442 365760 2858
rect 367066 2854 367094 3060
rect 368170 2938 368198 3060
rect 368170 2910 368336 2938
rect 367054 2848 367106 2854
rect 367054 2790 367106 2796
rect 368202 2816 368258 2825
rect 368202 2751 368258 2760
rect 366824 1556 366876 1562
rect 366824 1498 366876 1504
rect 365732 1414 365852 1442
rect 365824 480 365852 1414
rect 366836 762 366864 1498
rect 366836 734 367048 762
rect 367020 480 367048 734
rect 368216 480 368244 2751
rect 368308 1562 368336 2910
rect 369274 2825 369302 3060
rect 370056 2922 370176 2938
rect 370378 2922 370406 3060
rect 370044 2916 370176 2922
rect 370096 2910 370176 2916
rect 370044 2858 370096 2864
rect 369260 2816 369316 2825
rect 369260 2751 369316 2760
rect 369030 2680 369086 2689
rect 369086 2638 369440 2666
rect 369030 2615 369086 2624
rect 368296 1556 368348 1562
rect 368296 1498 368348 1504
rect 369412 480 369440 2638
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 2615
rect 380360 1562 380388 2774
rect 380912 1578 380940 2790
rect 381404 2751 381460 2760
rect 382292 1578 382320 2858
rect 383626 2802 383654 3060
rect 384730 2904 384758 3060
rect 385834 2922 385862 3060
rect 385822 2916 385874 2922
rect 384730 2876 384988 2904
rect 384960 2825 384988 2876
rect 385822 2858 385874 2864
rect 383476 2780 383528 2786
rect 383476 2722 383528 2728
rect 383580 2774 383654 2802
rect 384762 2816 384818 2825
rect 383488 1578 383516 2722
rect 383580 2553 383608 2774
rect 384762 2751 384818 2760
rect 384946 2816 385002 2825
rect 386938 2802 386966 3060
rect 388042 2825 388070 3060
rect 389146 2854 389174 3060
rect 389134 2848 389186 2854
rect 387154 2816 387210 2825
rect 386938 2774 387012 2802
rect 384946 2751 385002 2760
rect 383566 2544 383622 2553
rect 383566 2479 383622 2488
rect 380348 1556 380400 1562
rect 380912 1550 381216 1578
rect 382292 1550 382412 1578
rect 383488 1550 383608 1578
rect 380348 1498 380400 1504
rect 381188 480 381216 1550
rect 382384 480 382412 1550
rect 383580 480 383608 1550
rect 384776 480 384804 2751
rect 386984 1562 387012 2774
rect 387154 2751 387210 2760
rect 387798 2816 387854 2825
rect 387798 2751 387854 2760
rect 388028 2816 388084 2825
rect 389134 2790 389186 2796
rect 390250 2802 390278 3060
rect 391354 2961 391382 3060
rect 392458 2961 392486 3060
rect 391340 2952 391396 2961
rect 392444 2952 392500 2961
rect 391340 2887 391396 2896
rect 391848 2916 391900 2922
rect 393562 2938 393590 3060
rect 392444 2887 392500 2896
rect 393228 2916 393280 2922
rect 391848 2858 391900 2864
rect 393562 2910 393636 2938
rect 394666 2922 394694 3060
rect 393228 2858 393280 2864
rect 390250 2774 390324 2802
rect 388028 2751 388084 2760
rect 385776 1556 385828 1562
rect 385776 1498 385828 1504
rect 386972 1556 387024 1562
rect 386972 1498 387024 1504
rect 385788 762 385816 1498
rect 385788 734 386000 762
rect 385972 480 386000 734
rect 387168 480 387196 2751
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 2751
rect 389454 2544 389510 2553
rect 389454 2479 389510 2488
rect 389468 480 389496 2479
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390296 105 390324 2774
rect 390558 2680 390614 2689
rect 390614 2638 390692 2666
rect 390558 2615 390614 2624
rect 390664 480 390692 2638
rect 391860 480 391888 2858
rect 393240 2825 393268 2858
rect 393504 2848 393556 2854
rect 393226 2816 393282 2825
rect 393226 2751 393282 2760
rect 393502 2816 393504 2825
rect 393556 2816 393558 2825
rect 393502 2751 393558 2760
rect 393608 1562 393636 2910
rect 394056 2916 394108 2922
rect 394654 2916 394706 2922
rect 394108 2876 394280 2904
rect 394056 2858 394108 2864
rect 392676 1556 392728 1562
rect 392676 1498 392728 1504
rect 393596 1556 393648 1562
rect 393596 1498 393648 1504
rect 390282 96 390338 105
rect 390282 31 390338 40
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396170 96 396226 105
rect 396510 82 396622 480
rect 396226 54 396622 82
rect 396170 31 396226 40
rect 396510 -960 396622 54
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405660 377 405688 2774
rect 406810 2802 406838 3060
rect 407914 2802 407942 3060
rect 409018 2961 409046 3060
rect 409004 2952 409060 2961
rect 409004 2887 409060 2896
rect 410122 2825 410150 3060
rect 409602 2816 409658 2825
rect 406810 2774 406884 2802
rect 407914 2774 407988 2802
rect 406014 2751 406070 2760
rect 406028 480 406056 2751
rect 406856 1329 406884 2774
rect 406842 1320 406898 1329
rect 406842 1255 406898 1264
rect 407210 640 407266 649
rect 407210 575 407266 584
rect 407224 480 407252 575
rect 405646 368 405702 377
rect 405646 303 405702 312
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 407960 105 407988 2774
rect 409602 2751 409658 2760
rect 410108 2816 410164 2825
rect 411226 2802 411254 3060
rect 410108 2751 410164 2760
rect 411180 2774 411254 2802
rect 411720 2848 411772 2854
rect 411720 2790 411772 2796
rect 412330 2802 412358 3060
rect 413434 2802 413462 3060
rect 414538 2802 414566 3060
rect 415642 2802 415670 3060
rect 416594 2816 416650 2825
rect 408406 2000 408462 2009
rect 408406 1935 408462 1944
rect 408420 480 408448 1935
rect 409616 480 409644 2751
rect 410430 2680 410486 2689
rect 410486 2638 410840 2666
rect 410430 2615 410486 2624
rect 410812 480 410840 2638
rect 411180 649 411208 2774
rect 411732 1578 411760 2790
rect 412330 2774 412404 2802
rect 413434 2774 413508 2802
rect 414538 2774 414612 2802
rect 415642 2774 415716 2802
rect 411732 1550 411944 1578
rect 411166 640 411222 649
rect 411166 575 411222 584
rect 411916 480 411944 1550
rect 412376 921 412404 2774
rect 413480 1057 413508 2774
rect 414294 1320 414350 1329
rect 414294 1255 414350 1264
rect 413466 1048 413522 1057
rect 413466 983 413522 992
rect 412362 912 412418 921
rect 412362 847 412418 856
rect 414308 480 414336 1255
rect 414584 513 414612 2774
rect 415688 1329 415716 2774
rect 416746 2802 416774 3060
rect 416594 2751 416650 2760
rect 416700 2774 416774 2802
rect 417850 2802 417878 3060
rect 417974 2816 418030 2825
rect 417850 2774 417924 2802
rect 415674 1320 415730 1329
rect 415674 1255 415730 1264
rect 416608 1034 416636 2751
rect 416700 1193 416728 2774
rect 416686 1184 416742 1193
rect 416686 1119 416742 1128
rect 416608 1006 416728 1034
rect 414570 504 414626 513
rect 407946 96 408002 105
rect 407946 31 408002 40
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412822 368 412878 377
rect 413070 354 413182 480
rect 412878 326 413182 354
rect 412822 303 412878 312
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 416700 480 416728 1006
rect 417896 785 417924 2774
rect 418954 2802 418982 3060
rect 420058 2802 420086 3060
rect 421162 2961 421190 3060
rect 421148 2952 421204 2961
rect 421148 2887 421204 2896
rect 422266 2802 422294 3060
rect 423370 2825 423398 3060
rect 418954 2774 419028 2802
rect 420058 2774 420132 2802
rect 417974 2751 418030 2760
rect 417882 776 417938 785
rect 417882 711 417938 720
rect 417988 626 418016 2751
rect 419000 2009 419028 2774
rect 418986 2000 419042 2009
rect 418986 1935 419042 1944
rect 420104 649 420132 2774
rect 422220 2774 422294 2802
rect 423356 2816 423412 2825
rect 421378 1048 421434 1057
rect 421378 983 421434 992
rect 420182 912 420238 921
rect 420182 847 420238 856
rect 417896 598 418016 626
rect 418986 640 419042 649
rect 417896 480 417924 598
rect 418986 575 419042 584
rect 420090 640 420146 649
rect 420090 575 420146 584
rect 419000 480 419028 575
rect 420196 480 420224 847
rect 421392 480 421420 983
rect 414570 439 414626 448
rect 415306 96 415362 105
rect 415462 82 415574 480
rect 415362 54 415574 82
rect 415306 31 415362 40
rect 415462 -960 415574 54
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422220 134 422248 2774
rect 424474 2802 424502 3060
rect 425578 2802 425606 3060
rect 426682 2802 426710 3060
rect 427786 2802 427814 3060
rect 424474 2774 424548 2802
rect 425578 2774 425652 2802
rect 426682 2774 426756 2802
rect 423356 2751 423412 2760
rect 424520 2145 424548 2774
rect 424506 2136 424562 2145
rect 424506 2071 424562 2080
rect 425624 1329 425652 2774
rect 423770 1320 423826 1329
rect 423770 1255 423826 1264
rect 425610 1320 425666 1329
rect 425610 1255 425666 1264
rect 423784 480 423812 1255
rect 424966 1184 425022 1193
rect 424966 1119 425022 1128
rect 424980 480 425008 1119
rect 426162 776 426218 785
rect 426162 711 426218 720
rect 426176 480 426204 711
rect 422546 354 422658 480
rect 422758 368 422814 377
rect 422546 326 422758 354
rect 422208 128 422260 134
rect 422208 70 422260 76
rect 422546 -960 422658 326
rect 422758 303 422814 312
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426728 241 426756 2774
rect 427740 2774 427814 2802
rect 428890 2802 428918 3060
rect 429994 2802 430022 3060
rect 431098 2802 431126 3060
rect 432050 2816 432106 2825
rect 428890 2774 428964 2802
rect 429994 2774 430068 2802
rect 431098 2774 431172 2802
rect 427740 2009 427768 2774
rect 427266 2000 427322 2009
rect 427266 1935 427322 1944
rect 427726 2000 427782 2009
rect 427726 1935 427782 1944
rect 427280 480 427308 1935
rect 428462 640 428518 649
rect 428462 575 428518 584
rect 428476 480 428504 575
rect 426714 232 426770 241
rect 426714 167 426770 176
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435376 241 435404 598
rect 435560 480 435588 598
rect 436756 480 436784 1935
rect 435362 232 435418 241
rect 435362 167 435418 176
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437478 368 437534 377
rect 437910 354 438022 480
rect 437534 326 438022 354
rect 437478 303 437534 312
rect 437910 -960 438022 326
rect 438780 202 438808 2774
rect 439134 2544 439190 2553
rect 439134 2479 439190 2488
rect 439148 480 439176 2479
rect 439976 1873 440004 2774
rect 441080 2689 441108 2774
rect 441066 2680 441122 2689
rect 441066 2615 441122 2624
rect 442184 2553 442212 2774
rect 442170 2544 442226 2553
rect 442170 2479 442226 2488
rect 443288 2417 443316 2774
rect 444300 2774 444374 2802
rect 445450 2802 445478 3060
rect 446554 2802 446582 3060
rect 447658 2802 447686 3060
rect 448762 2802 448790 3060
rect 449866 2854 449894 3060
rect 449854 2848 449906 2854
rect 445450 2774 445524 2802
rect 446554 2774 446628 2802
rect 447658 2774 447732 2802
rect 448762 2774 448836 2802
rect 449854 2790 449906 2796
rect 450970 2802 450998 3060
rect 452074 2961 452102 3060
rect 453178 2961 453206 3060
rect 452060 2952 452116 2961
rect 452060 2887 452116 2896
rect 453164 2952 453220 2961
rect 453164 2887 453220 2896
rect 454282 2802 454310 3060
rect 455386 2961 455414 3060
rect 456490 2961 456518 3060
rect 455372 2952 455428 2961
rect 455372 2887 455428 2896
rect 456476 2952 456532 2961
rect 456476 2887 456532 2896
rect 450970 2774 451044 2802
rect 454282 2774 454356 2802
rect 442630 2408 442686 2417
rect 442630 2343 442686 2352
rect 443274 2408 443330 2417
rect 443274 2343 443330 2352
rect 439962 1864 440018 1873
rect 439962 1799 440018 1808
rect 439964 1352 440016 1358
rect 439964 1294 440016 1300
rect 438768 196 438820 202
rect 438768 138 438820 144
rect 439106 -960 439218 480
rect 439976 218 440004 1294
rect 441526 1184 441582 1193
rect 441526 1119 441582 1128
rect 441540 480 441568 1119
rect 442644 480 442672 2343
rect 443826 1728 443882 1737
rect 443826 1663 443882 1672
rect 443840 480 443868 1663
rect 440302 218 440414 480
rect 439976 190 440414 218
rect 440302 -960 440414 190
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444300 134 444328 2774
rect 445496 2281 445524 2774
rect 445022 2272 445078 2281
rect 445022 2207 445078 2216
rect 445482 2272 445538 2281
rect 445482 2207 445538 2216
rect 445036 480 445064 2207
rect 446600 2145 446628 2774
rect 446218 2136 446274 2145
rect 446218 2071 446274 2080
rect 446586 2136 446642 2145
rect 446586 2071 446642 2080
rect 446232 480 446260 2071
rect 447414 2000 447470 2009
rect 447414 1935 447470 1944
rect 447428 480 447456 1935
rect 447704 513 447732 2774
rect 448808 2009 448836 2774
rect 450910 2680 450966 2689
rect 450910 2615 450966 2624
rect 448794 2000 448850 2009
rect 448794 1935 448850 1944
rect 449806 1864 449862 1873
rect 449806 1799 449862 1808
rect 447690 504 447746 513
rect 444288 128 444340 134
rect 444288 70 444340 76
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 449820 480 449848 1799
rect 450924 480 450952 2615
rect 451016 1358 451044 2774
rect 452106 2544 452162 2553
rect 452106 2479 452162 2488
rect 451004 1352 451056 1358
rect 451004 1294 451056 1300
rect 452120 480 452148 2479
rect 453302 2408 453358 2417
rect 453302 2343 453358 2352
rect 453316 480 453344 2343
rect 454328 1290 454356 2774
rect 457594 2774 457622 3060
rect 458698 2961 458726 3060
rect 459802 2961 459830 3060
rect 458684 2952 458740 2961
rect 458684 2887 458740 2896
rect 459788 2952 459844 2961
rect 459788 2887 459844 2896
rect 460388 2848 460440 2854
rect 460388 2790 460440 2796
rect 457594 2746 457668 2774
rect 455694 2272 455750 2281
rect 455694 2207 455750 2216
rect 454316 1284 454368 1290
rect 454316 1226 454368 1232
rect 455708 480 455736 2207
rect 456890 2136 456946 2145
rect 456890 2071 456946 2080
rect 456904 480 456932 2071
rect 447690 439 447746 448
rect 448582 218 448694 480
rect 448440 202 448694 218
rect 448428 196 448694 202
rect 448480 190 448694 196
rect 448428 138 448480 144
rect 448582 -960 448694 190
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454132 128 454184 134
rect 454470 82 454582 480
rect 454184 76 454582 82
rect 454132 70 454582 76
rect 454144 54 454582 70
rect 454470 -960 454582 54
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457640 105 457668 2746
rect 459190 2000 459246 2009
rect 459190 1935 459246 1944
rect 457916 598 458128 626
rect 457718 504 457774 513
rect 457916 490 457944 598
rect 457774 462 457944 490
rect 458100 480 458128 598
rect 459204 480 459232 1935
rect 460400 480 460428 2790
rect 460906 2774 460934 3060
rect 460860 2746 460934 2774
rect 462010 2774 462038 3060
rect 463114 2774 463142 3060
rect 464218 2961 464246 3060
rect 464204 2952 464260 2961
rect 464204 2887 464260 2896
rect 463974 2816 464030 2825
rect 462010 2746 462084 2774
rect 463114 2746 463188 2774
rect 463974 2751 464030 2760
rect 465322 2774 465350 3060
rect 466426 2774 466454 3060
rect 467530 2802 467558 3060
rect 468634 2802 468662 3060
rect 469738 2802 469766 3060
rect 470842 2938 470870 3060
rect 471946 2961 471974 3060
rect 471932 2952 471988 2961
rect 470842 2910 471284 2938
rect 471256 2825 471284 2910
rect 471932 2887 471988 2896
rect 469862 2816 469918 2825
rect 467530 2774 467604 2802
rect 468634 2774 468708 2802
rect 469738 2774 469812 2802
rect 457718 439 457774 448
rect 457626 96 457682 105
rect 457626 31 457682 40
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 460860 134 460888 2746
rect 462056 1358 462084 2746
rect 462686 2680 462742 2689
rect 462742 2638 462820 2666
rect 462686 2615 462742 2624
rect 461308 1352 461360 1358
rect 461308 1294 461360 1300
rect 462044 1352 462096 1358
rect 462044 1294 462096 1300
rect 461320 762 461348 1294
rect 461320 734 461624 762
rect 461596 480 461624 734
rect 462792 480 462820 2638
rect 463160 2281 463188 2746
rect 463146 2272 463202 2281
rect 463146 2207 463202 2216
rect 463988 480 464016 2751
rect 465322 2746 465396 2774
rect 465080 1284 465132 1290
rect 465132 1244 465212 1272
rect 465080 1226 465132 1232
rect 465184 480 465212 1244
rect 465368 513 465396 2746
rect 466380 2746 466454 2774
rect 466274 2544 466330 2553
rect 466274 2479 466330 2488
rect 465354 504 465410 513
rect 460848 128 460900 134
rect 460848 70 460900 76
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466288 480 466316 2479
rect 466380 1222 466408 2746
rect 467286 2544 467342 2553
rect 467342 2502 467512 2530
rect 467286 2479 467342 2488
rect 466368 1216 466420 1222
rect 466368 1158 466420 1164
rect 467484 480 467512 2502
rect 467576 1358 467604 2774
rect 468680 2145 468708 2774
rect 468666 2136 468722 2145
rect 468666 2071 468722 2080
rect 469784 2009 469812 2774
rect 469862 2751 469918 2760
rect 471058 2816 471114 2825
rect 471058 2751 471114 2760
rect 471242 2816 471298 2825
rect 473050 2802 473078 3060
rect 474154 2802 474182 3060
rect 475258 2802 475286 3060
rect 476362 2802 476390 3060
rect 477466 2802 477494 3060
rect 473050 2774 473124 2802
rect 474154 2774 474228 2802
rect 475258 2774 475332 2802
rect 471242 2751 471298 2760
rect 469770 2000 469826 2009
rect 469770 1935 469826 1944
rect 467564 1352 467616 1358
rect 467564 1294 467616 1300
rect 468496 598 468708 626
rect 465354 439 465410 448
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468496 105 468524 598
rect 468680 480 468708 598
rect 469876 480 469904 2751
rect 471072 480 471100 2751
rect 473096 1358 473124 2774
rect 472992 1352 473044 1358
rect 472992 1294 473044 1300
rect 473084 1352 473136 1358
rect 473084 1294 473136 1300
rect 473004 1154 473032 1294
rect 473360 1284 473412 1290
rect 473360 1226 473412 1232
rect 472992 1148 473044 1154
rect 472992 1090 473044 1096
rect 473372 626 473400 1226
rect 473372 598 473492 626
rect 473464 480 473492 598
rect 468482 96 468538 105
rect 468482 31 468538 40
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 82 472338 480
rect 472440 128 472492 134
rect 472226 76 472440 82
rect 472226 70 472492 76
rect 472226 54 472480 70
rect 472226 -960 472338 54
rect 473422 -960 473534 480
rect 474200 202 474228 2774
rect 474554 2272 474610 2281
rect 474554 2207 474610 2216
rect 474568 480 474596 2207
rect 475304 785 475332 2774
rect 476316 2774 476390 2802
rect 477420 2774 477494 2802
rect 478570 2802 478598 3060
rect 478880 2848 478932 2854
rect 478570 2774 478644 2802
rect 478880 2790 478932 2796
rect 479674 2802 479702 3060
rect 480778 2802 480806 3060
rect 481882 2802 481910 3060
rect 482834 2816 482890 2825
rect 475382 2680 475438 2689
rect 475438 2638 475792 2666
rect 475382 2615 475438 2624
rect 475290 776 475346 785
rect 475290 711 475346 720
rect 475764 480 475792 2638
rect 474188 196 474240 202
rect 474188 138 474240 144
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476316 105 476344 2774
rect 476394 504 476450 513
rect 476450 462 476528 490
rect 476394 439 476450 448
rect 476500 354 476528 462
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476302 96 476358 105
rect 476302 31 476358 40
rect 476918 -960 477030 326
rect 477420 134 477448 2774
rect 477868 1216 477920 1222
rect 477868 1158 477920 1164
rect 477880 626 477908 1158
rect 477880 598 478184 626
rect 478156 480 478184 598
rect 478616 513 478644 2774
rect 478892 1358 478920 2790
rect 479674 2774 479748 2802
rect 480778 2774 480852 2802
rect 481882 2774 481956 2802
rect 479720 1358 479748 2774
rect 480534 2136 480590 2145
rect 480534 2071 480590 2080
rect 478880 1352 478932 1358
rect 478880 1294 478932 1300
rect 479708 1352 479760 1358
rect 479708 1294 479760 1300
rect 478892 1154 479012 1170
rect 478880 1148 479012 1154
rect 478932 1142 479012 1148
rect 478880 1090 478932 1096
rect 478602 504 478658 513
rect 477408 128 477460 134
rect 477408 70 477460 76
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484228 270 484256 2774
rect 485240 480 485268 2790
rect 486160 2774 486326 2802
rect 487264 2774 487430 2802
rect 488460 2774 488534 2802
rect 489610 2802 489638 3060
rect 490714 2802 490742 3060
rect 491818 2825 491846 3060
rect 489610 2774 489684 2802
rect 484216 264 484268 270
rect 484216 206 484268 212
rect 485198 -960 485310 480
rect 486160 377 486188 2774
rect 486146 368 486202 377
rect 486146 303 486202 312
rect 486394 218 486506 480
rect 487264 241 487292 2774
rect 488460 1290 488488 2774
rect 488448 1284 488500 1290
rect 488448 1226 488500 1232
rect 487618 776 487674 785
rect 487618 711 487674 720
rect 487632 480 487660 711
rect 487250 232 487306 241
rect 486394 202 486648 218
rect 486394 196 486660 202
rect 486394 190 486608 196
rect 486394 -960 486506 190
rect 487250 167 487306 176
rect 486608 138 486660 144
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 493980 134 494008 2774
rect 496280 1358 496308 2774
rect 496268 1352 496320 1358
rect 496268 1294 496320 1300
rect 494702 912 494758 921
rect 494702 847 494758 856
rect 494716 480 494744 847
rect 497384 746 497412 2774
rect 498198 2544 498254 2553
rect 498198 2479 498254 2488
rect 497372 740 497424 746
rect 497372 682 497424 688
rect 495900 672 495952 678
rect 495900 614 495952 620
rect 495912 480 495940 614
rect 498212 480 498240 2479
rect 498488 649 498516 2774
rect 499500 2774 499574 2802
rect 500650 2802 500678 3060
rect 501754 2802 501782 3060
rect 502858 2802 502886 3060
rect 503962 2802 503990 3060
rect 505066 2802 505094 3060
rect 500650 2774 500724 2802
rect 501754 2774 502104 2802
rect 499500 678 499528 2774
rect 500696 814 500724 2774
rect 501696 1284 501748 1290
rect 501696 1226 501748 1232
rect 500684 808 500736 814
rect 500684 750 500736 756
rect 499488 672 499540 678
rect 498474 640 498530 649
rect 501708 660 501736 1226
rect 501708 632 501828 660
rect 499488 614 499540 620
rect 498474 575 498530 584
rect 500328 598 500632 626
rect 493968 128 494020 134
rect 493968 70 494020 76
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 218 497178 480
rect 497280 264 497332 270
rect 497066 212 497280 218
rect 497066 206 497332 212
rect 497066 190 497320 206
rect 497066 -960 497178 190
rect 498170 -960 498282 480
rect 498934 368 498990 377
rect 499366 354 499478 480
rect 498990 326 499478 354
rect 498934 303 498990 312
rect 499366 -960 499478 326
rect 500328 241 500356 598
rect 500604 480 500632 598
rect 501800 480 501828 632
rect 500314 232 500370 241
rect 500314 167 500370 176
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502076 377 502104 2774
rect 502720 2774 502886 2802
rect 503732 2774 503990 2802
rect 505020 2774 505094 2802
rect 505374 2816 505430 2825
rect 502062 368 502118 377
rect 502062 303 502118 312
rect 502720 241 502748 2774
rect 502706 232 502762 241
rect 502706 167 502762 176
rect 502954 82 503066 480
rect 503732 105 503760 2774
rect 504150 218 504262 480
rect 505020 270 505048 2774
rect 506170 2802 506198 3060
rect 507274 2802 507302 3060
rect 508378 2961 508406 3060
rect 508364 2952 508420 2961
rect 508364 2887 508420 2896
rect 509482 2825 509510 3060
rect 506170 2774 506244 2802
rect 505374 2751 505430 2760
rect 505388 480 505416 2751
rect 503824 202 504262 218
rect 505008 264 505060 270
rect 505008 206 505060 212
rect 503812 196 504262 202
rect 503864 190 504262 196
rect 503812 138 503864 144
rect 503166 96 503222 105
rect 502954 54 503166 82
rect 502954 -960 503066 54
rect 503166 31 503222 40
rect 503718 96 503774 105
rect 503718 31 503774 40
rect 504150 -960 504262 190
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 1294
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 510540 134 510568 2774
rect 513898 2802 513926 3060
rect 515002 2961 515030 3060
rect 514988 2952 515044 2961
rect 514988 2887 515044 2896
rect 516106 2802 516134 3060
rect 513898 2774 513972 2802
rect 512780 2751 512836 2760
rect 513944 746 513972 2774
rect 516060 2774 516134 2802
rect 517210 2802 517238 3060
rect 518314 2961 518342 3060
rect 518300 2952 518356 2961
rect 518300 2887 518356 2896
rect 519418 2802 519446 3060
rect 517210 2774 517376 2802
rect 516060 1290 516088 2774
rect 516048 1284 516100 1290
rect 516048 1226 516100 1232
rect 514760 808 514812 814
rect 514760 750 514812 756
rect 513932 740 513984 746
rect 513932 682 513984 688
rect 512458 640 512514 649
rect 512458 575 512514 584
rect 512472 480 512500 575
rect 514772 480 514800 750
rect 517150 640 517206 649
rect 517150 575 517206 584
rect 517164 480 517192 575
rect 511234 354 511346 480
rect 511448 468 511500 474
rect 511448 410 511500 416
rect 511460 354 511488 410
rect 511234 326 511488 354
rect 510528 128 510580 134
rect 510528 70 510580 76
rect 511234 -960 511346 326
rect 512430 -960 512542 480
rect 513534 354 513646 480
rect 513392 338 513646 354
rect 513380 332 513646 338
rect 513432 326 513646 332
rect 513380 274 513432 280
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515494 368 515550 377
rect 515926 354 516038 480
rect 515550 326 516038 354
rect 515494 303 515550 312
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 218 521926 480
rect 521672 202 521926 218
rect 522776 202 522804 2774
rect 523038 2544 523094 2553
rect 523038 2479 523094 2488
rect 523052 480 523080 2479
rect 521660 196 521926 202
rect 521712 190 521926 196
rect 521660 138 521712 144
rect 521814 -960 521926 190
rect 522764 196 522816 202
rect 522764 138 522816 144
rect 523010 -960 523122 480
rect 523880 406 523908 2774
rect 524234 2751 524290 2760
rect 526042 2774 526070 3060
rect 527146 2774 527174 3060
rect 524248 480 524276 2751
rect 526042 2746 526116 2774
rect 523868 400 523920 406
rect 523868 342 523920 348
rect 524206 -960 524318 480
rect 525402 82 525514 480
rect 526088 241 526116 2746
rect 527100 2746 527174 2774
rect 528250 2774 528278 3060
rect 529354 2961 529382 3060
rect 529340 2952 529396 2961
rect 529340 2887 529396 2896
rect 530458 2774 530486 3060
rect 531562 2961 531590 3060
rect 531548 2952 531604 2961
rect 531548 2887 531604 2896
rect 532666 2774 532694 3060
rect 528250 2746 528324 2774
rect 530458 2746 530532 2774
rect 526534 2680 526590 2689
rect 526590 2638 526668 2666
rect 526534 2615 526590 2624
rect 526640 480 526668 2638
rect 526074 232 526130 241
rect 526074 167 526130 176
rect 525616 128 525668 134
rect 525402 76 525616 82
rect 525402 70 525668 76
rect 525402 54 525656 70
rect 525402 -960 525514 54
rect 526598 -960 526710 480
rect 527100 134 527128 2746
rect 527638 2680 527694 2689
rect 527694 2638 527864 2666
rect 527638 2615 527694 2624
rect 527836 480 527864 2638
rect 528296 2009 528324 2746
rect 530030 2680 530086 2689
rect 530086 2638 530164 2666
rect 530030 2615 530086 2624
rect 528282 2000 528338 2009
rect 528282 1935 528338 1944
rect 529020 740 529072 746
rect 529020 682 529072 688
rect 529032 480 529060 682
rect 530136 480 530164 2638
rect 530504 1222 530532 2746
rect 532620 2746 532694 2774
rect 533770 2774 533798 3060
rect 534874 2802 534902 3060
rect 535978 2961 536006 3060
rect 535964 2952 536020 2961
rect 535964 2887 536020 2896
rect 537082 2802 537110 3060
rect 538186 2802 538214 3060
rect 534874 2774 534948 2802
rect 537082 2774 537156 2802
rect 533770 2746 533844 2774
rect 531320 1284 531372 1290
rect 531320 1226 531372 1232
rect 530492 1216 530544 1222
rect 530492 1158 530544 1164
rect 531332 480 531360 1226
rect 532620 626 532648 2746
rect 533342 2680 533398 2689
rect 533398 2638 533752 2666
rect 533342 2615 533398 2624
rect 532620 598 532740 626
rect 527088 128 527140 134
rect 527088 70 527140 76
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 354 532598 480
rect 532160 338 532598 354
rect 532712 338 532740 598
rect 533724 480 533752 2638
rect 533816 1358 533844 2746
rect 533804 1352 533856 1358
rect 533804 1294 533856 1300
rect 534920 785 534948 2774
rect 537128 1290 537156 2774
rect 538140 2774 538214 2802
rect 539290 2802 539318 3060
rect 540394 2802 540422 3060
rect 541498 2961 541526 3060
rect 541484 2952 541540 2961
rect 541484 2887 541540 2896
rect 542602 2825 542630 3060
rect 540794 2816 540850 2825
rect 539290 2774 539364 2802
rect 540394 2774 540468 2802
rect 537116 1284 537168 1290
rect 537116 1226 537168 1232
rect 537036 1154 537248 1170
rect 537024 1148 537248 1154
rect 537076 1142 537248 1148
rect 537024 1090 537076 1096
rect 534906 776 534962 785
rect 534906 711 534962 720
rect 534736 598 534948 626
rect 532148 332 532598 338
rect 532200 326 532598 332
rect 532148 274 532200 280
rect 532486 -960 532598 326
rect 532700 332 532752 338
rect 532700 274 532752 280
rect 533682 -960 533794 480
rect 534736 105 534764 598
rect 534920 480 534948 598
rect 537220 480 537248 1142
rect 534722 96 534778 105
rect 534722 31 534778 40
rect 534878 -960 534990 480
rect 536074 218 536186 480
rect 536288 264 536340 270
rect 536074 212 536288 218
rect 536074 206 536340 212
rect 536074 190 536328 206
rect 536074 -960 536186 190
rect 537178 -960 537290 480
rect 538140 270 538168 2774
rect 538128 264 538180 270
rect 538374 218 538486 480
rect 539336 474 539364 2774
rect 539324 468 539376 474
rect 539324 410 539376 416
rect 538128 206 538180 212
rect 538232 202 538486 218
rect 538220 196 538486 202
rect 538272 190 538486 196
rect 538220 138 538272 144
rect 538374 -960 538486 190
rect 539570 354 539682 480
rect 539784 400 539836 406
rect 539570 348 539784 354
rect 539570 342 539836 348
rect 539570 326 539824 342
rect 539570 -960 539682 326
rect 540440 202 540468 2774
rect 540794 2751 540850 2760
rect 542588 2816 542644 2825
rect 543706 2802 543734 3060
rect 542588 2751 542644 2760
rect 543660 2774 543734 2802
rect 544810 2774 544838 3060
rect 545914 2774 545942 3060
rect 547018 2774 547046 3060
rect 548122 2961 548150 3060
rect 548108 2952 548164 2961
rect 548108 2887 548164 2896
rect 549226 2774 549254 3060
rect 540808 480 540836 2751
rect 540428 196 540480 202
rect 540428 138 540480 144
rect 540766 -960 540878 480
rect 541962 218 542074 480
rect 542174 232 542230 241
rect 541962 190 542174 218
rect 541962 -960 542074 190
rect 542174 167 542230 176
rect 542820 128 542872 134
rect 543158 82 543270 480
rect 543660 134 543688 2774
rect 544810 2746 544884 2774
rect 545914 2746 545988 2774
rect 547018 2746 547092 2774
rect 544382 2000 544438 2009
rect 544382 1935 544438 1944
rect 544396 480 544424 1935
rect 542872 76 543270 82
rect 542820 70 543270 76
rect 543648 128 543700 134
rect 543648 70 543700 76
rect 542832 54 543270 70
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 544856 105 544884 2746
rect 545302 2544 545358 2553
rect 545358 2502 545528 2530
rect 545302 2479 545358 2488
rect 545500 480 545528 2502
rect 545960 785 545988 2746
rect 546500 1216 546552 1222
rect 546500 1158 546552 1164
rect 545946 776 546002 785
rect 545946 711 546002 720
rect 544842 96 544898 105
rect 544842 31 544898 40
rect 545458 -960 545570 480
rect 546512 354 546540 1158
rect 546654 354 546766 480
rect 547064 406 547092 2746
rect 549180 2746 549254 2774
rect 550330 2774 550358 3060
rect 551434 2774 551462 3060
rect 550330 2746 550404 2774
rect 547878 2544 547934 2553
rect 547878 2479 547934 2488
rect 547892 480 547920 2479
rect 549180 1154 549208 2746
rect 550088 1352 550140 1358
rect 550088 1294 550140 1300
rect 549168 1148 549220 1154
rect 549168 1090 549220 1096
rect 550100 762 550128 1294
rect 550376 1290 550404 2746
rect 551388 2746 551462 2774
rect 552538 2774 552566 3060
rect 553642 2802 553670 3060
rect 554746 2802 554774 3060
rect 553642 2774 553716 2802
rect 552538 2746 552612 2774
rect 550364 1284 550416 1290
rect 550364 1226 550416 1232
rect 550100 734 550312 762
rect 550284 480 550312 734
rect 551388 649 551416 2746
rect 552478 2680 552534 2689
rect 552478 2615 552534 2624
rect 552492 762 552520 2615
rect 552584 921 552612 2746
rect 553688 1358 553716 2774
rect 554700 2774 554774 2802
rect 555850 2802 555878 3060
rect 556954 2802 556982 3060
rect 555850 2774 555924 2802
rect 553676 1352 553728 1358
rect 553676 1294 553728 1300
rect 553768 1216 553820 1222
rect 553768 1158 553820 1164
rect 552570 912 552626 921
rect 552570 847 552626 856
rect 552492 734 552704 762
rect 551374 640 551430 649
rect 551374 575 551430 584
rect 551480 598 551692 626
rect 551480 480 551508 598
rect 546512 326 546766 354
rect 547052 400 547104 406
rect 547052 342 547104 348
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 354 549158 480
rect 548720 338 549158 354
rect 548708 332 549158 338
rect 548760 326 549158 332
rect 548708 274 548760 280
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 551664 377 551692 598
rect 552676 480 552704 734
rect 553780 480 553808 1158
rect 551650 368 551706 377
rect 551650 303 551706 312
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554700 338 554728 2774
rect 555896 1222 555924 2774
rect 556908 2774 556982 2802
rect 558058 2802 558086 3060
rect 558550 2816 558606 2825
rect 558058 2774 558132 2802
rect 555884 1216 555936 1222
rect 555884 1158 555936 1164
rect 554688 332 554740 338
rect 554688 274 554740 280
rect 554780 264 554832 270
rect 554934 218 555046 480
rect 554832 212 555046 218
rect 554780 206 555046 212
rect 554792 190 555046 206
rect 554934 -960 555046 190
rect 556130 354 556242 480
rect 556344 468 556396 474
rect 556344 410 556396 416
rect 556356 354 556384 410
rect 556130 326 556384 354
rect 556130 -960 556242 326
rect 556908 270 556936 2774
rect 556896 264 556948 270
rect 557326 218 557438 480
rect 558104 377 558132 2774
rect 559162 2802 559190 3060
rect 560266 2802 560294 3060
rect 559162 2774 559236 2802
rect 558550 2751 558606 2760
rect 558564 480 558592 2751
rect 559208 513 559236 2774
rect 560220 2774 560294 2802
rect 561370 2802 561398 3060
rect 562474 2802 562502 3060
rect 563578 2802 563606 3060
rect 565634 2816 565690 2825
rect 561370 2774 561444 2802
rect 562474 2774 562548 2802
rect 563578 2774 563652 2802
rect 559286 2544 559342 2553
rect 559342 2502 559420 2530
rect 559286 2479 559342 2488
rect 559194 504 559250 513
rect 558090 368 558146 377
rect 558090 303 558146 312
rect 556896 206 556948 212
rect 557000 202 557438 218
rect 556988 196 557438 202
rect 557040 190 557438 196
rect 556988 138 557040 144
rect 557326 -960 557438 190
rect 558522 -960 558634 480
rect 559194 439 559250 448
rect 559392 354 559420 2502
rect 559718 354 559830 480
rect 559392 326 559830 354
rect 559718 -960 559830 326
rect 560220 202 560248 2774
rect 560208 196 560260 202
rect 560208 138 560260 144
rect 560484 128 560536 134
rect 560822 82 560934 480
rect 561416 134 561444 2774
rect 560536 76 560934 82
rect 560484 70 560934 76
rect 561404 128 561456 134
rect 561404 70 561456 76
rect 562018 82 562130 480
rect 562520 241 562548 2774
rect 563242 776 563298 785
rect 563242 711 563298 720
rect 563256 480 563284 711
rect 562506 232 562562 241
rect 562506 167 562562 176
rect 562230 96 562286 105
rect 560496 54 560934 70
rect 560822 -960 560934 54
rect 562018 54 562230 82
rect 562018 -960 562130 54
rect 562230 31 562286 40
rect 563214 -960 563326 480
rect 563624 105 563652 2774
rect 565634 2751 565690 2760
rect 565648 480 565676 2751
rect 571064 1352 571116 1358
rect 571064 1294 571116 1300
rect 567568 1284 567620 1290
rect 567568 1226 567620 1232
rect 566832 1148 566884 1154
rect 566832 1090 566884 1096
rect 566844 480 566872 1090
rect 564410 354 564522 480
rect 564624 400 564676 406
rect 564410 348 564624 354
rect 564410 342 564676 348
rect 564410 326 564664 342
rect 563610 96 563666 105
rect 563610 31 563666 40
rect 564410 -960 564522 326
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 1226
rect 570326 912 570382 921
rect 570326 847 570382 856
rect 569130 640 569186 649
rect 569130 575 569186 584
rect 569144 480 569172 575
rect 570340 480 570368 847
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571076 354 571104 1294
rect 573364 1216 573416 1222
rect 573364 1158 573416 1164
rect 571494 354 571606 480
rect 571076 326 571606 354
rect 571494 -960 571606 326
rect 572690 354 572802 480
rect 573376 354 573404 1158
rect 577134 504 577190 513
rect 573886 354 573998 480
rect 572690 338 572944 354
rect 572690 332 572956 338
rect 572690 326 572904 332
rect 572690 -960 572802 326
rect 573376 326 573998 354
rect 572904 274 572956 280
rect 573886 -960 573998 326
rect 575082 218 575194 480
rect 575754 368 575810 377
rect 576278 354 576390 480
rect 577134 439 577190 448
rect 575810 326 576390 354
rect 577148 354 577176 439
rect 577382 354 577494 480
rect 577148 326 577494 354
rect 575754 303 575810 312
rect 575296 264 575348 270
rect 575082 212 575296 218
rect 575082 206 575348 212
rect 575082 190 575336 206
rect 575082 -960 575194 190
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 218 578690 480
rect 578578 202 578832 218
rect 578578 196 578844 202
rect 578578 190 578792 196
rect 578578 -960 578690 190
rect 578792 138 578844 144
rect 579774 -960 579886 480
rect 580970 82 581082 480
rect 581826 232 581882 241
rect 582166 218 582278 480
rect 581882 190 582278 218
rect 581826 167 581882 176
rect 581184 128 581236 134
rect 580970 76 581184 82
rect 580970 70 581236 76
rect 580970 54 581224 70
rect 580970 -960 581082 54
rect 582166 -960 582278 190
rect 583362 82 583474 480
rect 583574 96 583630 105
rect 583362 54 583574 82
rect 583362 -960 583474 54
rect 583574 31 583630 40
<< via2 >>
rect 85486 680040 85542 680096
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 250442 680312 250498 680368
rect 241426 679496 241482 679552
rect 72606 623464 72662 623520
rect 3514 619112 3570 619168
rect 3422 606056 3478 606112
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 72790 615168 72846 615224
rect 72882 611088 72938 611144
rect 74446 627680 74502 627736
rect 73066 619384 73122 619440
rect 72974 606872 73030 606928
rect 232778 623464 232834 623520
rect 232318 619384 232374 619440
rect 232686 619384 232742 619440
rect 233146 627680 233202 627736
rect 232870 615168 232926 615224
rect 232962 611088 233018 611144
rect 235262 627952 235318 628008
rect 232410 606872 232466 606928
rect 233054 606872 233110 606928
rect 72698 602792 72754 602848
rect 233146 602792 233202 602848
rect 72974 598576 73030 598632
rect 231766 598576 231822 598632
rect 72882 594496 72938 594552
rect 72698 586200 72754 586256
rect 71778 577904 71834 577960
rect 73066 590280 73122 590336
rect 73066 581984 73122 582040
rect 233054 594496 233110 594552
rect 232778 590280 232834 590336
rect 232870 586200 232926 586256
rect 75826 577516 75882 577552
rect 75826 577496 75828 577516
rect 75828 577496 75880 577516
rect 75880 577496 75882 577516
rect 3606 514800 3662 514856
rect 3514 501744 3570 501800
rect 3514 462576 3570 462632
rect 3514 449520 3570 449576
rect 3146 410488 3202 410544
rect 3606 409400 3662 409456
rect 3514 409264 3570 409320
rect 3422 405864 3478 405920
rect 3606 406000 3662 406056
rect 3514 397432 3570 397488
rect 17130 359216 17186 359272
rect 3606 358400 3662 358456
rect 3422 345344 3478 345400
rect 17038 332288 17094 332344
rect 17038 330384 17094 330440
rect 3422 321000 3478 321056
rect 3330 149776 3386 149832
rect 3238 97552 3294 97608
rect 3790 320864 3846 320920
rect 3606 320728 3662 320784
rect 3514 293120 3570 293176
rect 3514 289040 3570 289096
rect 3790 306176 3846 306232
rect 3606 254088 3662 254144
rect 3514 241032 3570 241088
rect 3514 201864 3570 201920
rect 17222 358264 17278 358320
rect 17774 356088 17830 356144
rect 17682 355136 17738 355192
rect 17498 353368 17554 353424
rect 17406 352280 17462 352336
rect 16854 240896 16910 240952
rect 16762 239944 16818 240000
rect 16946 213968 17002 214024
rect 16946 212064 17002 212120
rect 17590 350512 17646 350568
rect 17498 235048 17554 235104
rect 17406 233960 17462 234016
rect 72790 409128 72846 409184
rect 71686 407804 71688 407824
rect 71688 407804 71740 407824
rect 71740 407804 71742 407824
rect 71686 407768 71742 407804
rect 66166 407632 66222 407688
rect 64510 407224 64566 407280
rect 140686 407940 140688 407960
rect 140688 407940 140740 407960
rect 140740 407940 140742 407960
rect 140686 407904 140742 407940
rect 52366 407108 52422 407144
rect 52366 407088 52368 407108
rect 52368 407088 52420 407108
rect 52420 407088 52422 407108
rect 56506 407088 56562 407144
rect 59266 407088 59322 407144
rect 99286 407088 99342 407144
rect 108946 407088 109002 407144
rect 111706 407088 111762 407144
rect 114466 407088 114522 407144
rect 117226 407088 117282 407144
rect 118606 407088 118662 407144
rect 121366 407088 121422 407144
rect 124126 407088 124182 407144
rect 126886 407088 126942 407144
rect 139306 407088 139362 407144
rect 151358 407124 151360 407144
rect 151360 407124 151412 407144
rect 151412 407124 151414 407144
rect 151358 407088 151414 407124
rect 86222 406580 86224 406600
rect 86224 406580 86276 406600
rect 86276 406580 86278 406600
rect 86222 406544 86278 406580
rect 88614 406544 88670 406600
rect 95974 406544 96030 406600
rect 81070 406428 81126 406464
rect 81070 406408 81072 406428
rect 81072 406408 81124 406428
rect 81124 406408 81126 406428
rect 83646 406408 83702 406464
rect 48686 406136 48742 406192
rect 53470 406136 53526 406192
rect 61106 406136 61162 406192
rect 17866 330656 17922 330712
rect 17774 237768 17830 237824
rect 17682 236816 17738 236872
rect 17590 232192 17646 232248
rect 143354 321952 143410 322008
rect 19430 321136 19486 321192
rect 17866 212336 17922 212392
rect 3514 188808 3570 188864
rect 3606 136720 3662 136776
rect 3514 84632 3570 84688
rect 3422 58520 3478 58576
rect 3606 45464 3662 45520
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 18694 319640 18750 319696
rect 19430 316104 19486 316160
rect 19798 316240 19854 316296
rect 19798 315832 19854 315888
rect 19798 306584 19854 306640
rect 19798 306176 19854 306232
rect 19798 296928 19854 296984
rect 19798 296520 19854 296576
rect 19706 209616 19762 209672
rect 19706 209344 19762 209400
rect 62762 321564 62818 321600
rect 62762 321544 62764 321564
rect 62764 321544 62816 321564
rect 62816 321544 62818 321564
rect 63866 321544 63922 321600
rect 67638 321544 67694 321600
rect 44178 320084 44180 320104
rect 44180 320084 44232 320104
rect 44232 320084 44234 320104
rect 44178 320048 44234 320084
rect 45006 320048 45062 320104
rect 50158 320068 50214 320104
rect 50158 320048 50160 320068
rect 50160 320048 50212 320068
rect 50212 320048 50214 320068
rect 36082 319912 36138 319968
rect 39578 319912 39634 319968
rect 36542 319096 36598 319152
rect 37922 319096 37978 319152
rect 40682 319252 40738 319288
rect 40682 319232 40684 319252
rect 40684 319232 40736 319252
rect 40736 319232 40738 319252
rect 42062 319232 42118 319288
rect 51262 320068 51318 320104
rect 51262 320048 51264 320068
rect 51264 320048 51316 320068
rect 51316 320048 51318 320068
rect 52366 320048 52422 320104
rect 53470 320048 53526 320104
rect 56506 319640 56562 319696
rect 59358 320048 59414 320104
rect 60646 320048 60702 320104
rect 67638 320456 67694 320512
rect 65338 320048 65394 320104
rect 68650 320048 68706 320104
rect 71134 320048 71190 320104
rect 59910 319912 59966 319968
rect 60830 319912 60886 319968
rect 66442 319912 66498 319968
rect 70398 319232 70454 319288
rect 46202 319096 46258 319152
rect 46202 318824 46258 318880
rect 48318 291080 48374 291136
rect 52366 291080 52422 291136
rect 53746 291080 53802 291136
rect 56506 291080 56562 291136
rect 59266 291080 59322 291136
rect 62026 291080 62082 291136
rect 64786 291080 64842 291136
rect 68926 291080 68982 291136
rect 66166 290672 66222 290728
rect 74630 320456 74686 320512
rect 72146 320048 72202 320104
rect 73342 320048 73398 320104
rect 75734 320048 75790 320104
rect 71686 291080 71742 291136
rect 73986 290264 74042 290320
rect 79230 320084 79232 320104
rect 79232 320084 79284 320104
rect 79284 320084 79286 320104
rect 79230 320048 79286 320084
rect 78678 319640 78734 319696
rect 77298 319232 77354 319288
rect 77206 291080 77262 291136
rect 78586 291080 78642 291136
rect 81346 291080 81402 291136
rect 84106 291080 84162 291136
rect 86866 291080 86922 291136
rect 89626 291080 89682 291136
rect 91006 291080 91062 291136
rect 93766 291080 93822 291136
rect 99286 291080 99342 291136
rect 106186 291116 106188 291136
rect 106188 291116 106240 291136
rect 106240 291116 106242 291136
rect 106186 291080 106242 291116
rect 102046 290944 102102 291000
rect 143262 320456 143318 320512
rect 157338 318960 157394 319016
rect 117226 291080 117282 291136
rect 114466 290944 114522 291000
rect 111706 290844 111708 290864
rect 111708 290844 111760 290864
rect 111760 290844 111762 290864
rect 111706 290808 111762 290844
rect 140686 290808 140742 290864
rect 104806 290672 104862 290728
rect 118606 290672 118662 290728
rect 121366 290264 121422 290320
rect 96526 290128 96582 290184
rect 126886 290400 126942 290456
rect 139306 290400 139362 290456
rect 108946 289992 109002 290048
rect 122838 289992 122894 290048
rect 46202 287680 46258 287736
rect 150898 287408 150954 287464
rect 142066 203768 142122 203824
rect 69754 203496 69810 203552
rect 71134 203496 71190 203552
rect 72238 203496 72294 203552
rect 73342 203496 73398 203552
rect 74354 203496 74410 203552
rect 75734 203496 75790 203552
rect 78034 203496 78090 203552
rect 76930 202972 76986 203008
rect 76930 202952 76932 202972
rect 76932 202952 76984 202972
rect 76984 202952 76986 202972
rect 41602 202136 41658 202192
rect 35898 201320 35954 201376
rect 36542 201340 36598 201376
rect 36542 201320 36544 201340
rect 36544 201320 36596 201340
rect 36596 201320 36598 201340
rect 37278 201356 37280 201376
rect 37280 201356 37332 201376
rect 37332 201356 37334 201376
rect 37278 201320 37334 201356
rect 38658 201320 38714 201376
rect 40038 201320 40094 201376
rect 44178 201320 44234 201376
rect 44362 201320 44418 201376
rect 63498 201320 63554 201376
rect 67638 201320 67694 201376
rect 79966 201320 80022 201376
rect 51078 201184 51134 201240
rect 52458 201184 52514 201240
rect 55586 201184 55642 201240
rect 59358 201184 59414 201240
rect 62118 201204 62174 201240
rect 62118 201184 62120 201204
rect 62120 201184 62172 201204
rect 62172 201184 62174 201204
rect 59450 201068 59506 201104
rect 59450 201048 59452 201068
rect 59452 201048 59504 201068
rect 59504 201048 59506 201068
rect 49698 200776 49754 200832
rect 51170 200796 51226 200832
rect 51170 200776 51172 200796
rect 51172 200776 51224 200796
rect 51224 200776 51226 200796
rect 62026 200640 62082 200696
rect 66258 200368 66314 200424
rect 64878 200252 64934 200288
rect 64878 200232 64880 200252
rect 64880 200232 64932 200252
rect 64932 200232 64934 200252
rect 213826 408448 213882 408504
rect 216586 408448 216642 408504
rect 233054 581984 233110 582040
rect 233146 577904 233202 577960
rect 235262 577516 235318 577552
rect 235262 577496 235264 577516
rect 235264 577496 235316 577516
rect 235316 577496 235318 577516
rect 226246 408448 226302 408504
rect 228822 408448 228878 408504
rect 222106 408312 222162 408368
rect 223486 408312 223542 408368
rect 159362 401648 159418 401704
rect 159086 341672 159142 341728
rect 158718 340040 158774 340096
rect 158810 338680 158866 338736
rect 158718 221720 158774 221776
rect 158994 337184 159050 337240
rect 158902 335960 158958 336016
rect 158810 220380 158866 220416
rect 158810 220360 158812 220380
rect 158812 220360 158864 220380
rect 158864 220360 158866 220380
rect 209502 407088 209558 407144
rect 211066 407088 211122 407144
rect 218978 407088 219034 407144
rect 231766 407088 231822 407144
rect 234526 407088 234582 407144
rect 237286 407088 237342 407144
rect 177210 359216 177266 359272
rect 176658 330792 176714 330848
rect 177118 330384 177174 330440
rect 160006 283192 160062 283248
rect 159086 223352 159142 223408
rect 159362 223352 159418 223408
rect 158994 218864 159050 218920
rect 158902 217640 158958 217696
rect 158902 216688 158958 216744
rect 159454 221720 159510 221776
rect 159546 216688 159602 216744
rect 142066 201184 142122 201240
rect 143446 201184 143502 201240
rect 143446 200796 143502 200832
rect 143446 200776 143448 200796
rect 143448 200776 143500 200796
rect 143500 200776 143502 200796
rect 177394 358264 177450 358320
rect 177854 356088 177910 356144
rect 177762 355136 177818 355192
rect 177670 353368 177726 353424
rect 177578 352280 177634 352336
rect 177486 350512 177542 350568
rect 177210 240896 177266 240952
rect 177394 253816 177450 253872
rect 177394 244024 177450 244080
rect 177302 239944 177358 240000
rect 177394 237768 177450 237824
rect 177118 232192 177174 232248
rect 177026 212336 177082 212392
rect 177486 236816 177542 236872
rect 177946 332288 178002 332344
rect 177946 330384 178002 330440
rect 178130 321272 178186 321328
rect 178038 320592 178094 320648
rect 177762 244232 177818 244288
rect 177670 235048 177726 235104
rect 177578 233960 177634 234016
rect 177762 234640 177818 234696
rect 177762 232192 177818 232248
rect 177854 213968 177910 214024
rect 177854 212064 177910 212120
rect 178038 319368 178094 319424
rect 238574 406544 238630 406600
rect 241426 407088 241482 407144
rect 251086 408448 251142 408504
rect 253846 408448 253902 408504
rect 259366 408448 259422 408504
rect 264886 408448 264942 408504
rect 266266 408448 266322 408504
rect 274546 408448 274602 408504
rect 271786 408312 271842 408368
rect 269026 408040 269082 408096
rect 246946 407088 247002 407144
rect 249706 407088 249762 407144
rect 256606 407088 256662 407144
rect 262126 407088 262182 407144
rect 243726 406544 243782 406600
rect 276846 407088 276902 407144
rect 278686 408448 278742 408504
rect 281078 406544 281134 406600
rect 284206 407088 284262 407144
rect 286506 408312 286562 408368
rect 299386 407124 299388 407144
rect 299388 407124 299440 407144
rect 299440 407124 299442 407144
rect 299386 407088 299442 407124
rect 300766 407088 300822 407144
rect 318062 407768 318118 407824
rect 317418 407088 317474 407144
rect 316866 406000 316922 406056
rect 223486 321952 223542 322008
rect 228638 321952 228694 322008
rect 179786 321816 179842 321872
rect 179418 321716 179420 321736
rect 179420 321716 179472 321736
rect 179472 321716 179474 321736
rect 179418 321680 179474 321716
rect 226338 321716 226340 321736
rect 226340 321716 226392 321736
rect 226392 321716 226394 321736
rect 226338 321680 226394 321716
rect 179510 321544 179566 321600
rect 178958 321408 179014 321464
rect 178590 320184 178646 320240
rect 178774 320184 178830 320240
rect 178682 267688 178738 267744
rect 178406 205808 178462 205864
rect 178682 205808 178738 205864
rect 179510 321136 179566 321192
rect 179510 320184 179566 320240
rect 179326 205808 179382 205864
rect 179326 203768 179382 203824
rect 179602 243888 179658 243944
rect 179602 236408 179658 236464
rect 180154 321408 180210 321464
rect 200762 320084 200764 320104
rect 200764 320084 200816 320104
rect 200816 320084 200818 320104
rect 200762 320048 200818 320084
rect 196070 319368 196126 319424
rect 197358 319368 197414 319424
rect 198738 319368 198794 319424
rect 180522 318824 180578 318880
rect 195978 318860 195980 318880
rect 195980 318860 196032 318880
rect 196032 318860 196034 318880
rect 195978 318824 196034 318860
rect 201498 319232 201554 319288
rect 219438 321428 219494 321464
rect 219438 321408 219440 321428
rect 219440 321408 219492 321428
rect 219492 321408 219494 321428
rect 220450 321408 220506 321464
rect 207294 320592 207350 320648
rect 203154 320048 203210 320104
rect 203798 320048 203854 320104
rect 204350 320048 204406 320104
rect 204258 319096 204314 319152
rect 180338 287428 180394 287464
rect 211802 320048 211858 320104
rect 210422 319796 210478 319832
rect 210422 319776 210424 319796
rect 210424 319776 210476 319796
rect 210476 319776 210478 319796
rect 206282 319232 206338 319288
rect 209042 319232 209098 319288
rect 209318 291080 209374 291136
rect 211342 319116 211398 319152
rect 211342 319096 211344 319116
rect 211344 319096 211396 319116
rect 211396 319096 211398 319116
rect 211066 291080 211122 291136
rect 215114 319912 215170 319968
rect 213182 319368 213238 319424
rect 211986 319096 212042 319152
rect 213826 291080 213882 291136
rect 216402 319640 216458 319696
rect 216678 319640 216734 319696
rect 217874 319640 217930 319696
rect 218058 319640 218114 319696
rect 219254 319640 219310 319696
rect 216494 291080 216550 291136
rect 221830 320592 221886 320648
rect 224130 320084 224132 320104
rect 224132 320084 224184 320104
rect 224184 320084 224186 320104
rect 224130 320048 224186 320084
rect 227534 320048 227590 320104
rect 222842 319368 222898 319424
rect 219346 291080 219402 291136
rect 222106 291080 222162 291136
rect 226982 319912 227038 319968
rect 225602 319232 225658 319288
rect 223486 291080 223542 291136
rect 226246 291080 226302 291136
rect 228914 291080 228970 291136
rect 231214 320048 231270 320104
rect 229558 319932 229614 319968
rect 229558 319912 229560 319932
rect 229560 319912 229612 319932
rect 229612 319912 229614 319932
rect 231858 319660 231914 319696
rect 231858 319640 231860 319660
rect 231860 319640 231912 319660
rect 231912 319640 231914 319660
rect 232502 319640 232558 319696
rect 231766 291080 231822 291136
rect 236642 319504 236698 319560
rect 234066 319232 234122 319288
rect 235262 319268 235264 319288
rect 235264 319268 235316 319288
rect 235316 319268 235318 319288
rect 235262 319232 235318 319268
rect 233882 318824 233938 318880
rect 238022 319096 238078 319152
rect 239402 318960 239458 319016
rect 238666 291080 238722 291136
rect 241426 291080 241482 291136
rect 244186 291080 244242 291136
rect 246946 291080 247002 291136
rect 249706 291080 249762 291136
rect 251086 291080 251142 291136
rect 253846 291080 253902 291136
rect 256606 291080 256662 291136
rect 259366 291080 259422 291136
rect 237286 290944 237342 291000
rect 264886 291080 264942 291136
rect 269026 291080 269082 291136
rect 271786 291080 271842 291136
rect 274546 291080 274602 291136
rect 277306 291080 277362 291136
rect 303066 319368 303122 319424
rect 302882 319232 302938 319288
rect 281446 291080 281502 291136
rect 284206 291080 284262 291136
rect 266266 290672 266322 290728
rect 278686 290672 278742 290728
rect 262126 290400 262182 290456
rect 234526 289992 234582 290048
rect 286598 289856 286654 289912
rect 299018 289856 299074 289912
rect 299662 289856 299718 289912
rect 310794 289856 310850 289912
rect 180338 287408 180340 287428
rect 180340 287408 180392 287428
rect 180392 287408 180394 287428
rect 229742 203496 229798 203552
rect 231122 203496 231178 203552
rect 232226 203496 232282 203552
rect 233330 203496 233386 203552
rect 234434 203496 234490 203552
rect 235722 203496 235778 203552
rect 237010 203496 237066 203552
rect 238022 203496 238078 203552
rect 318154 405864 318210 405920
rect 320086 401668 320142 401704
rect 320086 401648 320088 401668
rect 320088 401648 320140 401668
rect 320140 401648 320142 401668
rect 319534 341672 319590 341728
rect 319442 283192 319498 283248
rect 317418 223352 317474 223408
rect 317510 221720 317566 221776
rect 317602 217640 317658 217696
rect 195978 201320 196034 201376
rect 196162 201320 196218 201376
rect 197358 201320 197414 201376
rect 198738 201320 198794 201376
rect 200118 201320 200174 201376
rect 204350 201320 204406 201376
rect 211250 201320 211306 201376
rect 219990 201320 220046 201376
rect 222198 201340 222254 201376
rect 222198 201320 222200 201340
rect 222200 201320 222252 201340
rect 222252 201320 222254 201340
rect 178958 200368 179014 200424
rect 204258 201184 204314 201240
rect 211158 201048 211214 201104
rect 215298 201184 215354 201240
rect 219438 201184 219494 201240
rect 223578 201356 223580 201376
rect 223580 201356 223632 201376
rect 223632 201356 223634 201376
rect 223578 201320 223634 201356
rect 224958 201320 225014 201376
rect 238942 201320 238998 201376
rect 303158 201356 303160 201376
rect 303160 201356 303212 201376
rect 303212 201356 303214 201376
rect 303158 201320 303214 201356
rect 303526 201340 303582 201376
rect 303526 201320 303528 201340
rect 303528 201320 303580 201340
rect 303580 201320 303582 201340
rect 209870 200776 209926 200832
rect 201314 200504 201370 200560
rect 201498 200504 201554 200560
rect 201866 200504 201922 200560
rect 220818 200232 220874 200288
rect 201130 200096 201186 200152
rect 201314 200096 201370 200152
rect 318798 220768 318854 220824
rect 318798 220360 318854 220416
rect 318890 218864 318946 218920
rect 318890 218048 318946 218104
rect 319626 340040 319682 340096
rect 319718 338680 319774 338736
rect 319810 337184 319866 337240
rect 319902 335960 319958 336016
rect 319626 221720 319682 221776
rect 319718 220768 319774 220824
rect 319902 223352 319958 223408
rect 319810 218048 319866 218104
rect 319442 217640 319498 217696
rect 321098 406272 321154 406328
rect 321190 321000 321246 321056
rect 322754 409400 322810 409456
rect 322478 320864 322534 320920
rect 324962 289040 325018 289096
rect 325238 406408 325294 406464
rect 328090 320728 328146 320784
rect 329378 407632 329434 407688
rect 330942 409264 330998 409320
rect 330666 406136 330722 406192
rect 333334 408176 333390 408232
rect 334806 407224 334862 407280
rect 335082 407496 335138 407552
rect 336002 396208 336058 396264
rect 336094 380840 336150 380896
rect 336094 357040 336150 357096
rect 336370 407360 336426 407416
rect 336462 371184 336518 371240
rect 336370 355136 336426 355192
rect 336370 348064 336426 348120
rect 336278 341672 336334 341728
rect 336186 339768 336242 339824
rect 336186 331472 336242 331528
rect 336922 381520 336978 381576
rect 336922 379616 336978 379672
rect 337290 377576 337346 377632
rect 337106 376352 337162 376408
rect 336922 372544 336978 372600
rect 337290 369280 337346 369336
rect 336554 366696 336610 366752
rect 337290 366016 337346 366072
rect 337106 362208 337162 362264
rect 336922 360304 336978 360360
rect 336922 357720 336978 357776
rect 336922 353232 336978 353288
rect 337290 352028 337346 352064
rect 337290 352008 337292 352028
rect 337292 352008 337344 352028
rect 337344 352008 337346 352028
rect 336922 340992 336978 341048
rect 337290 340448 337346 340504
rect 337290 339088 337346 339144
rect 336738 338544 336794 338600
rect 337106 327528 337162 327584
rect 336922 320456 336978 320512
rect 336922 318552 336978 318608
rect 337106 310256 337162 310312
rect 337106 308896 337162 308952
rect 337658 397568 337714 397624
rect 337658 396888 337714 396944
rect 337750 395664 337806 395720
rect 337658 394984 337714 395040
rect 337750 394304 337806 394360
rect 337658 393624 337714 393680
rect 337750 393080 337806 393136
rect 337658 392400 337714 392456
rect 337658 391720 337714 391776
rect 337750 391176 337806 391232
rect 337658 390496 337714 390552
rect 337750 389816 337806 389872
rect 337658 389172 337660 389192
rect 337660 389172 337712 389192
rect 337712 389172 337714 389192
rect 337658 389136 337714 389172
rect 337750 388592 337806 388648
rect 337842 387912 337898 387968
rect 337658 387232 337714 387288
rect 337750 386688 337806 386744
rect 337658 386008 337714 386064
rect 337750 385328 337806 385384
rect 337658 384648 337714 384704
rect 337750 384104 337806 384160
rect 337658 383424 337714 383480
rect 337750 382744 337806 382800
rect 337658 382100 337660 382120
rect 337660 382100 337712 382120
rect 337712 382100 337714 382120
rect 337658 382064 337714 382100
rect 337750 380160 337806 380216
rect 337658 378936 337714 378992
rect 337750 378256 337806 378312
rect 337750 377032 337806 377088
rect 337658 375672 337714 375728
rect 337750 375128 337806 375184
rect 337658 374448 337714 374504
rect 337750 373768 337806 373824
rect 337658 373088 337714 373144
rect 337566 371864 337622 371920
rect 337658 370640 337714 370696
rect 337658 369960 337714 370016
rect 337658 368600 337714 368656
rect 337750 368056 337806 368112
rect 337750 367376 337806 367432
rect 337658 365472 337714 365528
rect 337750 364792 337806 364848
rect 337658 364112 337714 364168
rect 337750 363568 337806 363624
rect 337658 362908 337714 362944
rect 337658 362888 337660 362908
rect 337660 362888 337712 362908
rect 337712 362888 337714 362908
rect 337566 361528 337622 361584
rect 337658 360984 337714 361040
rect 337658 359624 337714 359680
rect 337474 359080 337530 359136
rect 337750 358400 337806 358456
rect 337658 356496 337714 356552
rect 337658 355816 337714 355872
rect 337750 354592 337806 354648
rect 337566 353912 337622 353968
rect 337474 346840 337530 346896
rect 337658 352552 337714 352608
rect 337658 351328 337714 351384
rect 337658 350648 337714 350704
rect 337750 349968 337806 350024
rect 337658 349424 337714 349480
rect 337750 348744 337806 348800
rect 337658 347520 337714 347576
rect 337658 346160 337714 346216
rect 337658 345480 337714 345536
rect 337750 344972 337752 344992
rect 337752 344972 337804 344992
rect 337804 344972 337806 344992
rect 337750 344936 337806 344972
rect 337658 344256 337714 344312
rect 337750 343576 337806 343632
rect 337658 343032 337714 343088
rect 337566 342352 337622 342408
rect 337750 337864 337806 337920
rect 337658 337184 337714 337240
rect 337842 336504 337898 336560
rect 337658 335960 337714 336016
rect 337566 335280 337622 335336
rect 337750 334600 337806 334656
rect 337658 333920 337714 333976
rect 337750 333376 337806 333432
rect 337750 332696 337806 332752
rect 337658 332016 337714 332072
rect 337658 330792 337714 330848
rect 337750 330112 337806 330168
rect 337658 329432 337714 329488
rect 337658 328888 337714 328944
rect 337566 328208 337622 328264
rect 337658 327020 337660 327040
rect 337660 327020 337712 327040
rect 337712 327020 337714 327040
rect 337658 326984 337714 327020
rect 337658 326304 337714 326360
rect 337566 325624 337622 325680
rect 337658 324944 337714 325000
rect 337750 324400 337806 324456
rect 337658 323720 337714 323776
rect 337474 323040 337530 323096
rect 337750 322496 337806 322552
rect 337658 321816 337714 321872
rect 337658 321136 337714 321192
rect 337750 319912 337806 319968
rect 337658 319232 337714 319288
rect 337658 317872 337714 317928
rect 337566 317328 337622 317384
rect 337658 316648 337714 316704
rect 337750 315968 337806 316024
rect 337658 315424 337714 315480
rect 337658 314764 337714 314800
rect 337658 314744 337660 314764
rect 337660 314744 337712 314764
rect 337712 314744 337714 314764
rect 337658 314064 337714 314120
rect 337658 313384 337714 313440
rect 337750 312840 337806 312896
rect 337750 312160 337806 312216
rect 337658 311480 337714 311536
rect 337658 310936 337714 310992
rect 337658 309576 337714 309632
rect 337658 308352 337714 308408
rect 337382 307672 337438 307728
rect 337658 306992 337714 307048
rect 337750 306448 337806 306504
rect 337658 305768 337714 305824
rect 337750 305088 337806 305144
rect 337658 304408 337714 304464
rect 337750 303864 337806 303920
rect 337658 303184 337714 303240
rect 336922 302504 336978 302560
rect 337658 301824 337714 301880
rect 337474 301280 337530 301336
rect 337658 300600 337714 300656
rect 337382 299920 337438 299976
rect 337106 299376 337162 299432
rect 337290 298696 337346 298752
rect 337750 298016 337806 298072
rect 337658 297336 337714 297392
rect 336922 296792 336978 296848
rect 337658 296112 337714 296168
rect 337106 295432 337162 295488
rect 336922 294888 336978 294944
rect 337658 294208 337714 294264
rect 337658 293528 337714 293584
rect 337750 292848 337806 292904
rect 337658 292304 337714 292360
rect 337750 291624 337806 291680
rect 337474 290944 337530 291000
rect 337106 290400 337162 290456
rect 337658 289740 337714 289776
rect 337658 289720 337660 289740
rect 337660 289720 337712 289740
rect 337712 289720 337714 289740
rect 336922 287136 336978 287192
rect 336738 286456 336794 286512
rect 336278 280744 336334 280800
rect 336830 280064 336886 280120
rect 336738 279384 336794 279440
rect 337106 286728 337162 286784
rect 337290 285232 337346 285288
rect 337750 289040 337806 289096
rect 337658 288360 337714 288416
rect 337750 287816 337806 287872
rect 337474 286864 337530 286920
rect 337474 285776 337530 285832
rect 337014 277480 337070 277536
rect 337198 277480 337254 277536
rect 336186 270408 336242 270464
rect 337014 277344 337070 277400
rect 337106 274352 337162 274408
rect 337290 277344 337346 277400
rect 337290 277208 337346 277264
rect 337198 272992 337254 273048
rect 337106 271788 337162 271824
rect 337106 271768 337108 271788
rect 337108 271768 337160 271788
rect 337160 271768 337162 271788
rect 337014 269184 337070 269240
rect 337382 276256 337438 276312
rect 337382 274896 337438 274952
rect 337290 268504 337346 268560
rect 337474 265240 337530 265296
rect 337658 284552 337714 284608
rect 337658 283872 337714 283928
rect 337750 283328 337806 283384
rect 337658 282648 337714 282704
rect 337750 281968 337806 282024
rect 337658 281288 337714 281344
rect 337750 278840 337806 278896
rect 337658 278160 337714 278216
rect 337750 277480 337806 277536
rect 337842 277344 337898 277400
rect 337842 276800 337898 276856
rect 337842 275576 337898 275632
rect 337842 273672 337898 273728
rect 337842 272312 337898 272368
rect 337842 271088 337898 271144
rect 337842 269728 337898 269784
rect 338026 267824 338082 267880
rect 337934 267280 337990 267336
rect 337750 266600 337806 266656
rect 337658 265920 337714 265976
rect 337566 264696 337622 264752
rect 336830 264016 336886 264072
rect 337474 263336 337530 263392
rect 337382 262792 337438 262848
rect 337474 262112 337530 262168
rect 337658 261432 337714 261488
rect 337750 260752 337806 260808
rect 337658 260208 337714 260264
rect 337106 259528 337162 259584
rect 337658 258304 337714 258360
rect 339038 258576 339094 258632
rect 460018 409128 460074 409184
rect 472622 627680 472678 627736
rect 472530 623464 472586 623520
rect 472622 619384 472678 619440
rect 472530 615168 472586 615224
rect 472622 611088 472678 611144
rect 472438 606872 472494 606928
rect 472622 602792 472678 602848
rect 472622 590280 472678 590336
rect 472622 586200 472678 586256
rect 472622 577904 472678 577960
rect 472990 598576 473046 598632
rect 473082 594496 473138 594552
rect 473174 581984 473230 582040
rect 483478 680584 483534 680640
rect 510894 679156 510950 679212
rect 482006 381520 482062 381576
rect 482282 376896 482338 376952
rect 482374 367512 482430 367568
rect 482282 339632 482338 339688
rect 482466 362888 482522 362944
rect 482558 358264 482614 358320
rect 482650 353640 482706 353696
rect 482742 348880 482798 348936
rect 482926 395528 482982 395584
rect 580170 697176 580226 697232
rect 482926 390904 482982 390960
rect 580170 683848 580226 683904
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 482926 386316 482928 386336
rect 482928 386316 482980 386336
rect 482980 386316 482982 386336
rect 482926 386280 482982 386316
rect 580262 590960 580318 591016
rect 580170 577632 580226 577688
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 378392 580226 378448
rect 482926 372272 482982 372328
rect 580170 365064 580226 365120
rect 482834 344256 482890 344312
rect 482374 334872 482430 334928
rect 482282 330248 482338 330304
rect 482374 325624 482430 325680
rect 482282 320864 482338 320920
rect 482006 316240 482062 316296
rect 481914 264988 481970 265024
rect 481914 264968 481916 264988
rect 481916 264968 481968 264988
rect 481968 264968 481970 264988
rect 482098 311616 482154 311672
rect 352562 200640 352618 200696
rect 482190 306992 482246 307048
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 482926 302232 482982 302288
rect 482834 297608 482890 297664
rect 482742 292984 482798 293040
rect 482650 288224 482706 288280
rect 482558 283600 482614 283656
rect 482466 278976 482522 279032
rect 482374 274216 482430 274272
rect 482374 269592 482430 269648
rect 482282 260344 482338 260400
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 483473 680642 483539 680645
rect 483473 680640 486894 680642
rect 483473 680584 483478 680640
rect 483534 680584 486894 680640
rect 483473 680582 486894 680584
rect 483473 680579 483539 680582
rect 486834 680570 486894 680582
rect 250437 680370 250503 680373
rect 247940 680368 250503 680370
rect 247940 680312 250442 680368
rect 250498 680312 250503 680368
rect 247940 680310 250503 680312
rect 250437 680307 250503 680310
rect 85481 680098 85547 680101
rect 85376 680096 85547 680098
rect 85376 680040 85486 680096
rect 85542 680040 85547 680096
rect 85376 680038 85547 680040
rect 85481 680035 85547 680038
rect 240550 679554 240610 680068
rect 241421 679554 241487 679557
rect 240550 679552 241487 679554
rect 240550 679496 241426 679552
rect 241482 679496 241487 679552
rect 240550 679494 241487 679496
rect 241421 679491 241487 679494
rect 510889 679214 510955 679217
rect 510784 679212 510955 679214
rect 510784 679156 510894 679212
rect 510950 679156 510955 679212
rect 510784 679154 510955 679156
rect 510889 679151 510955 679154
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 235257 628010 235323 628013
rect 235214 628008 235323 628010
rect 235214 627952 235262 628008
rect 235318 627952 235323 628008
rect 235214 627947 235323 627952
rect 74441 627738 74507 627741
rect 233141 627738 233207 627741
rect 235214 627738 235274 627947
rect 74441 627736 75348 627738
rect 74441 627680 74446 627736
rect 74502 627680 75348 627736
rect 74441 627678 75348 627680
rect 233141 627736 235274 627738
rect 233141 627680 233146 627736
rect 233202 627708 235274 627736
rect 472617 627738 472683 627741
rect 472617 627736 474812 627738
rect 233202 627680 235244 627708
rect 233141 627678 235244 627680
rect 472617 627680 472622 627736
rect 472678 627680 474812 627736
rect 472617 627678 474812 627680
rect 74441 627675 74507 627678
rect 233141 627675 233207 627678
rect 472617 627675 472683 627678
rect 72601 623522 72667 623525
rect 232773 623522 232839 623525
rect 472525 623522 472591 623525
rect 72601 623520 75348 623522
rect 72601 623464 72606 623520
rect 72662 623464 75348 623520
rect 72601 623462 75348 623464
rect 232773 623520 235244 623522
rect 232773 623464 232778 623520
rect 232834 623464 235244 623520
rect 232773 623462 235244 623464
rect 472525 623520 474812 623522
rect 472525 623464 472530 623520
rect 472586 623464 474812 623520
rect 472525 623462 474812 623464
rect 72601 623459 72667 623462
rect 232773 623459 232839 623462
rect 472525 623459 472591 623462
rect 73061 619442 73127 619445
rect 232313 619442 232379 619445
rect 232681 619442 232747 619445
rect 472617 619442 472683 619445
rect 73061 619440 75348 619442
rect 73061 619384 73066 619440
rect 73122 619384 75348 619440
rect 73061 619382 75348 619384
rect 232313 619440 235244 619442
rect 232313 619384 232318 619440
rect 232374 619384 232686 619440
rect 232742 619384 235244 619440
rect 232313 619382 235244 619384
rect 472617 619440 474812 619442
rect 472617 619384 472622 619440
rect 472678 619384 474812 619440
rect 472617 619382 474812 619384
rect 73061 619379 73127 619382
rect 232313 619379 232379 619382
rect 232681 619379 232747 619382
rect 472617 619379 472683 619382
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 583520 617388 584960 617628
rect 72785 615226 72851 615229
rect 232865 615226 232931 615229
rect 472525 615226 472591 615229
rect 72785 615224 75348 615226
rect 72785 615168 72790 615224
rect 72846 615168 75348 615224
rect 72785 615166 75348 615168
rect 232865 615224 235244 615226
rect 232865 615168 232870 615224
rect 232926 615168 235244 615224
rect 232865 615166 235244 615168
rect 472525 615224 474812 615226
rect 472525 615168 472530 615224
rect 472586 615168 474812 615224
rect 472525 615166 474812 615168
rect 72785 615163 72851 615166
rect 232865 615163 232931 615166
rect 472525 615163 472591 615166
rect 72877 611146 72943 611149
rect 232957 611146 233023 611149
rect 472617 611146 472683 611149
rect 72877 611144 75348 611146
rect 72877 611088 72882 611144
rect 72938 611088 75348 611144
rect 72877 611086 75348 611088
rect 232957 611144 235244 611146
rect 232957 611088 232962 611144
rect 233018 611088 235244 611144
rect 232957 611086 235244 611088
rect 472617 611144 474812 611146
rect 472617 611088 472622 611144
rect 472678 611088 474812 611144
rect 472617 611086 474812 611088
rect 72877 611083 72943 611086
rect 232957 611083 233023 611086
rect 472617 611083 472683 611086
rect 72969 606930 73035 606933
rect 232405 606930 232471 606933
rect 233049 606930 233115 606933
rect 472433 606930 472499 606933
rect 72969 606928 75348 606930
rect 72969 606872 72974 606928
rect 73030 606872 75348 606928
rect 72969 606870 75348 606872
rect 232405 606928 235244 606930
rect 232405 606872 232410 606928
rect 232466 606872 233054 606928
rect 233110 606872 235244 606928
rect 232405 606870 235244 606872
rect 472433 606928 474812 606930
rect 472433 606872 472438 606928
rect 472494 606872 474812 606928
rect 472433 606870 474812 606872
rect 72969 606867 73035 606870
rect 232405 606867 232471 606870
rect 233049 606867 233115 606870
rect 472433 606867 472499 606870
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect 72693 602850 72759 602853
rect 233141 602850 233207 602853
rect 472617 602850 472683 602853
rect 72693 602848 75348 602850
rect 72693 602792 72698 602848
rect 72754 602792 75348 602848
rect 72693 602790 75348 602792
rect 233141 602848 235244 602850
rect 233141 602792 233146 602848
rect 233202 602792 235244 602848
rect 233141 602790 235244 602792
rect 472617 602848 474812 602850
rect 472617 602792 472622 602848
rect 472678 602792 474812 602848
rect 472617 602790 474812 602792
rect 72693 602787 72759 602790
rect 233141 602787 233207 602790
rect 472617 602787 472683 602790
rect 72969 598634 73035 598637
rect 231761 598634 231827 598637
rect 472985 598634 473051 598637
rect 72969 598632 75348 598634
rect 72969 598576 72974 598632
rect 73030 598576 75348 598632
rect 72969 598574 75348 598576
rect 231761 598632 235244 598634
rect 231761 598576 231766 598632
rect 231822 598576 235244 598632
rect 231761 598574 235244 598576
rect 472985 598632 474812 598634
rect 472985 598576 472990 598632
rect 473046 598576 474812 598632
rect 472985 598574 474812 598576
rect 72969 598571 73035 598574
rect 231761 598571 231827 598574
rect 472985 598571 473051 598574
rect 72877 594554 72943 594557
rect 233049 594554 233115 594557
rect 473077 594554 473143 594557
rect 72877 594552 75348 594554
rect 72877 594496 72882 594552
rect 72938 594496 75348 594552
rect 72877 594494 75348 594496
rect 233049 594552 235244 594554
rect 233049 594496 233054 594552
rect 233110 594496 235244 594552
rect 233049 594494 235244 594496
rect 473077 594552 474812 594554
rect 473077 594496 473082 594552
rect 473138 594496 474812 594552
rect 473077 594494 474812 594496
rect 72877 594491 72943 594494
rect 233049 594491 233115 594494
rect 473077 594491 473143 594494
rect -960 592908 480 593148
rect 580257 591018 580323 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 583520 590868 584960 590958
rect 73061 590338 73127 590341
rect 232773 590338 232839 590341
rect 472617 590338 472683 590341
rect 73061 590336 75348 590338
rect 73061 590280 73066 590336
rect 73122 590280 75348 590336
rect 73061 590278 75348 590280
rect 232773 590336 235244 590338
rect 232773 590280 232778 590336
rect 232834 590280 235244 590336
rect 232773 590278 235244 590280
rect 472617 590336 474812 590338
rect 472617 590280 472622 590336
rect 472678 590280 474812 590336
rect 472617 590278 474812 590280
rect 73061 590275 73127 590278
rect 232773 590275 232839 590278
rect 472617 590275 472683 590278
rect 72693 586258 72759 586261
rect 232865 586258 232931 586261
rect 472617 586258 472683 586261
rect 72693 586256 75348 586258
rect 72693 586200 72698 586256
rect 72754 586200 75348 586256
rect 72693 586198 75348 586200
rect 232865 586256 235244 586258
rect 232865 586200 232870 586256
rect 232926 586200 235244 586256
rect 232865 586198 235244 586200
rect 472617 586256 474812 586258
rect 472617 586200 472622 586256
rect 472678 586200 474812 586256
rect 472617 586198 474812 586200
rect 72693 586195 72759 586198
rect 232865 586195 232931 586198
rect 472617 586195 472683 586198
rect 73061 582042 73127 582045
rect 233049 582042 233115 582045
rect 473169 582042 473235 582045
rect 73061 582040 75348 582042
rect 73061 581984 73066 582040
rect 73122 581984 75348 582040
rect 73061 581982 75348 581984
rect 233049 582040 235244 582042
rect 233049 581984 233054 582040
rect 233110 581984 235244 582040
rect 233049 581982 235244 581984
rect 473169 582040 474812 582042
rect 473169 581984 473174 582040
rect 473230 581984 474812 582040
rect 473169 581982 474812 581984
rect 73061 581979 73127 581982
rect 233049 581979 233115 581982
rect 473169 581979 473235 581982
rect -960 579852 480 580092
rect 71773 577962 71839 577965
rect 233141 577962 233207 577965
rect 472617 577962 472683 577965
rect 71773 577960 75900 577962
rect 71773 577904 71778 577960
rect 71834 577932 75900 577960
rect 233141 577960 235244 577962
rect 71834 577904 75930 577932
rect 71773 577902 75930 577904
rect 71773 577899 71839 577902
rect 75870 577557 75930 577902
rect 233141 577904 233146 577960
rect 233202 577932 235244 577960
rect 472617 577960 474812 577962
rect 233202 577904 235274 577932
rect 233141 577902 235274 577904
rect 233141 577899 233207 577902
rect 75821 577552 75930 577557
rect 75821 577496 75826 577552
rect 75882 577496 75930 577552
rect 75821 577494 75930 577496
rect 235214 577557 235274 577902
rect 472617 577904 472622 577960
rect 472678 577904 474812 577960
rect 472617 577902 474812 577904
rect 472617 577899 472683 577902
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 235214 577552 235323 577557
rect 235214 577496 235262 577552
rect 235318 577496 235323 577552
rect 583520 577540 584960 577630
rect 235214 577494 235323 577496
rect 75821 577491 75887 577494
rect 235257 577491 235323 577494
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 583520 511172 584960 511412
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 3601 409458 3667 409461
rect 322749 409458 322815 409461
rect 3601 409456 322815 409458
rect 3601 409400 3606 409456
rect 3662 409400 322754 409456
rect 322810 409400 322815 409456
rect 3601 409398 322815 409400
rect 3601 409395 3667 409398
rect 322749 409395 322815 409398
rect 3509 409322 3575 409325
rect 330937 409322 331003 409325
rect 3509 409320 331003 409322
rect 3509 409264 3514 409320
rect 3570 409264 330942 409320
rect 330998 409264 331003 409320
rect 3509 409262 331003 409264
rect 3509 409259 3575 409262
rect 330937 409259 331003 409262
rect 72785 409186 72851 409189
rect 460013 409186 460079 409189
rect 72785 409184 460079 409186
rect 72785 409128 72790 409184
rect 72846 409128 460018 409184
rect 460074 409128 460079 409184
rect 72785 409126 460079 409128
rect 72785 409123 72851 409126
rect 460013 409123 460079 409126
rect 213494 408444 213500 408508
rect 213564 408506 213570 408508
rect 213821 408506 213887 408509
rect 213564 408504 213887 408506
rect 213564 408448 213826 408504
rect 213882 408448 213887 408504
rect 213564 408446 213887 408448
rect 213564 408444 213570 408446
rect 213821 408443 213887 408446
rect 216254 408444 216260 408508
rect 216324 408506 216330 408508
rect 216581 408506 216647 408509
rect 226241 408508 226307 408509
rect 216324 408504 216647 408506
rect 216324 408448 216586 408504
rect 216642 408448 216647 408504
rect 216324 408446 216647 408448
rect 216324 408444 216330 408446
rect 216581 408443 216647 408446
rect 226190 408444 226196 408508
rect 226260 408506 226307 408508
rect 226260 408504 226352 408506
rect 226302 408448 226352 408504
rect 226260 408446 226352 408448
rect 226260 408444 226307 408446
rect 228582 408444 228588 408508
rect 228652 408506 228658 408508
rect 228817 408506 228883 408509
rect 251081 408508 251147 408509
rect 228652 408504 228883 408506
rect 228652 408448 228822 408504
rect 228878 408448 228883 408504
rect 228652 408446 228883 408448
rect 228652 408444 228658 408446
rect 226241 408443 226307 408444
rect 228817 408443 228883 408446
rect 251030 408444 251036 408508
rect 251100 408506 251147 408508
rect 251100 408504 251192 408506
rect 251142 408448 251192 408504
rect 251100 408446 251192 408448
rect 251100 408444 251147 408446
rect 253606 408444 253612 408508
rect 253676 408506 253682 408508
rect 253841 408506 253907 408509
rect 253676 408504 253907 408506
rect 253676 408448 253846 408504
rect 253902 408448 253907 408504
rect 253676 408446 253907 408448
rect 253676 408444 253682 408446
rect 251081 408443 251147 408444
rect 253841 408443 253907 408446
rect 258574 408444 258580 408508
rect 258644 408506 258650 408508
rect 259361 408506 259427 408509
rect 258644 408504 259427 408506
rect 258644 408448 259366 408504
rect 259422 408448 259427 408504
rect 258644 408446 259427 408448
rect 258644 408444 258650 408446
rect 259361 408443 259427 408446
rect 263542 408444 263548 408508
rect 263612 408506 263618 408508
rect 264881 408506 264947 408509
rect 263612 408504 264947 408506
rect 263612 408448 264886 408504
rect 264942 408448 264947 408504
rect 263612 408446 264947 408448
rect 263612 408444 263618 408446
rect 264881 408443 264947 408446
rect 265934 408444 265940 408508
rect 266004 408506 266010 408508
rect 266261 408506 266327 408509
rect 266004 408504 266327 408506
rect 266004 408448 266266 408504
rect 266322 408448 266327 408504
rect 266004 408446 266327 408448
rect 266004 408444 266010 408446
rect 266261 408443 266327 408446
rect 273662 408444 273668 408508
rect 273732 408506 273738 408508
rect 274541 408506 274607 408509
rect 273732 408504 274607 408506
rect 273732 408448 274546 408504
rect 274602 408448 274607 408504
rect 273732 408446 274607 408448
rect 273732 408444 273738 408446
rect 274541 408443 274607 408446
rect 278446 408444 278452 408508
rect 278516 408506 278522 408508
rect 278681 408506 278747 408509
rect 278516 408504 278747 408506
rect 278516 408448 278686 408504
rect 278742 408448 278747 408504
rect 278516 408446 278747 408448
rect 278516 408444 278522 408446
rect 278681 408443 278747 408446
rect 221038 408308 221044 408372
rect 221108 408370 221114 408372
rect 222101 408370 222167 408373
rect 223481 408372 223547 408373
rect 221108 408368 222167 408370
rect 221108 408312 222106 408368
rect 222162 408312 222167 408368
rect 221108 408310 222167 408312
rect 221108 408308 221114 408310
rect 222101 408307 222167 408310
rect 223430 408308 223436 408372
rect 223500 408370 223547 408372
rect 223500 408368 223592 408370
rect 223542 408312 223592 408368
rect 223500 408310 223592 408312
rect 223500 408308 223547 408310
rect 271086 408308 271092 408372
rect 271156 408370 271162 408372
rect 271781 408370 271847 408373
rect 271156 408368 271847 408370
rect 271156 408312 271786 408368
rect 271842 408312 271847 408368
rect 271156 408310 271847 408312
rect 271156 408308 271162 408310
rect 223481 408307 223547 408308
rect 271781 408307 271847 408310
rect 286174 408308 286180 408372
rect 286244 408370 286250 408372
rect 286501 408370 286567 408373
rect 286244 408368 286567 408370
rect 286244 408312 286506 408368
rect 286562 408312 286567 408368
rect 286244 408310 286567 408312
rect 286244 408308 286250 408310
rect 286501 408307 286567 408310
rect 90950 408172 90956 408236
rect 91020 408234 91026 408236
rect 333329 408234 333395 408237
rect 91020 408232 333395 408234
rect 91020 408176 333334 408232
rect 333390 408176 333395 408232
rect 91020 408174 333395 408176
rect 91020 408172 91026 408174
rect 333329 408171 333395 408174
rect 268510 408036 268516 408100
rect 268580 408098 268586 408100
rect 269021 408098 269087 408101
rect 268580 408096 269087 408098
rect 268580 408040 269026 408096
rect 269082 408040 269087 408096
rect 268580 408038 269087 408040
rect 268580 408036 268586 408038
rect 269021 408035 269087 408038
rect 139710 407900 139716 407964
rect 139780 407962 139786 407964
rect 140681 407962 140747 407965
rect 139780 407960 140747 407962
rect 139780 407904 140686 407960
rect 140742 407904 140747 407960
rect 139780 407902 140747 407904
rect 139780 407900 139786 407902
rect 140681 407899 140747 407902
rect 71078 407764 71084 407828
rect 71148 407826 71154 407828
rect 71681 407826 71747 407829
rect 71148 407824 71747 407826
rect 71148 407768 71686 407824
rect 71742 407768 71747 407824
rect 71148 407766 71747 407768
rect 71148 407764 71154 407766
rect 71681 407763 71747 407766
rect 93526 407764 93532 407828
rect 93596 407826 93602 407828
rect 318057 407826 318123 407829
rect 93596 407824 318123 407826
rect 93596 407768 318062 407824
rect 318118 407768 318123 407824
rect 93596 407766 318123 407768
rect 93596 407764 93602 407766
rect 318057 407763 318123 407766
rect 66161 407692 66227 407693
rect 66110 407628 66116 407692
rect 66180 407690 66227 407692
rect 66180 407688 66272 407690
rect 66222 407632 66272 407688
rect 66180 407630 66272 407632
rect 66180 407628 66227 407630
rect 101070 407628 101076 407692
rect 101140 407690 101146 407692
rect 329373 407690 329439 407693
rect 101140 407688 329439 407690
rect 101140 407632 329378 407688
rect 329434 407632 329439 407688
rect 101140 407630 329439 407632
rect 101140 407628 101146 407630
rect 66161 407627 66227 407628
rect 329373 407627 329439 407630
rect 106038 407492 106044 407556
rect 106108 407554 106114 407556
rect 335077 407554 335143 407557
rect 106108 407552 335143 407554
rect 106108 407496 335082 407552
rect 335138 407496 335143 407552
rect 106108 407494 335143 407496
rect 106108 407492 106114 407494
rect 335077 407491 335143 407494
rect 103646 407356 103652 407420
rect 103716 407418 103722 407420
rect 336365 407418 336431 407421
rect 103716 407416 336431 407418
rect 103716 407360 336370 407416
rect 336426 407360 336431 407416
rect 103716 407358 336431 407360
rect 103716 407356 103722 407358
rect 336365 407355 336431 407358
rect 63534 407220 63540 407284
rect 63604 407282 63610 407284
rect 64505 407282 64571 407285
rect 63604 407280 64571 407282
rect 63604 407224 64510 407280
rect 64566 407224 64571 407280
rect 63604 407222 64571 407224
rect 63604 407220 63610 407222
rect 64505 407219 64571 407222
rect 68502 407220 68508 407284
rect 68572 407282 68578 407284
rect 334801 407282 334867 407285
rect 68572 407280 334867 407282
rect 68572 407224 334806 407280
rect 334862 407224 334867 407280
rect 68572 407222 334867 407224
rect 68572 407220 68578 407222
rect 334801 407219 334867 407222
rect 51022 407084 51028 407148
rect 51092 407146 51098 407148
rect 52361 407146 52427 407149
rect 51092 407144 52427 407146
rect 51092 407088 52366 407144
rect 52422 407088 52427 407144
rect 51092 407086 52427 407088
rect 51092 407084 51098 407086
rect 52361 407083 52427 407086
rect 56174 407084 56180 407148
rect 56244 407146 56250 407148
rect 56501 407146 56567 407149
rect 56244 407144 56567 407146
rect 56244 407088 56506 407144
rect 56562 407088 56567 407144
rect 56244 407086 56567 407088
rect 56244 407084 56250 407086
rect 56501 407083 56567 407086
rect 58566 407084 58572 407148
rect 58636 407146 58642 407148
rect 59261 407146 59327 407149
rect 58636 407144 59327 407146
rect 58636 407088 59266 407144
rect 59322 407088 59327 407144
rect 58636 407086 59327 407088
rect 58636 407084 58642 407086
rect 59261 407083 59327 407086
rect 98678 407084 98684 407148
rect 98748 407146 98754 407148
rect 99281 407146 99347 407149
rect 98748 407144 99347 407146
rect 98748 407088 99286 407144
rect 99342 407088 99347 407144
rect 98748 407086 99347 407088
rect 98748 407084 98754 407086
rect 99281 407083 99347 407086
rect 108430 407084 108436 407148
rect 108500 407146 108506 407148
rect 108941 407146 109007 407149
rect 108500 407144 109007 407146
rect 108500 407088 108946 407144
rect 109002 407088 109007 407144
rect 108500 407086 109007 407088
rect 108500 407084 108506 407086
rect 108941 407083 109007 407086
rect 111006 407084 111012 407148
rect 111076 407146 111082 407148
rect 111701 407146 111767 407149
rect 111076 407144 111767 407146
rect 111076 407088 111706 407144
rect 111762 407088 111767 407144
rect 111076 407086 111767 407088
rect 111076 407084 111082 407086
rect 111701 407083 111767 407086
rect 113582 407084 113588 407148
rect 113652 407146 113658 407148
rect 114461 407146 114527 407149
rect 113652 407144 114527 407146
rect 113652 407088 114466 407144
rect 114522 407088 114527 407144
rect 113652 407086 114527 407088
rect 113652 407084 113658 407086
rect 114461 407083 114527 407086
rect 115974 407084 115980 407148
rect 116044 407146 116050 407148
rect 117221 407146 117287 407149
rect 118601 407148 118667 407149
rect 116044 407144 117287 407146
rect 116044 407088 117226 407144
rect 117282 407088 117287 407144
rect 116044 407086 117287 407088
rect 116044 407084 116050 407086
rect 117221 407083 117287 407086
rect 118550 407084 118556 407148
rect 118620 407146 118667 407148
rect 118620 407144 118712 407146
rect 118662 407088 118712 407144
rect 118620 407086 118712 407088
rect 118620 407084 118667 407086
rect 121126 407084 121132 407148
rect 121196 407146 121202 407148
rect 121361 407146 121427 407149
rect 121196 407144 121427 407146
rect 121196 407088 121366 407144
rect 121422 407088 121427 407144
rect 121196 407086 121427 407088
rect 121196 407084 121202 407086
rect 118601 407083 118667 407084
rect 121361 407083 121427 407086
rect 123334 407084 123340 407148
rect 123404 407146 123410 407148
rect 124121 407146 124187 407149
rect 123404 407144 124187 407146
rect 123404 407088 124126 407144
rect 124182 407088 124187 407144
rect 123404 407086 124187 407088
rect 123404 407084 123410 407086
rect 124121 407083 124187 407086
rect 126094 407084 126100 407148
rect 126164 407146 126170 407148
rect 126881 407146 126947 407149
rect 126164 407144 126947 407146
rect 126164 407088 126886 407144
rect 126942 407088 126947 407144
rect 126164 407086 126947 407088
rect 126164 407084 126170 407086
rect 126881 407083 126947 407086
rect 138422 407084 138428 407148
rect 138492 407146 138498 407148
rect 139301 407146 139367 407149
rect 138492 407144 139367 407146
rect 138492 407088 139306 407144
rect 139362 407088 139367 407144
rect 138492 407086 139367 407088
rect 138492 407084 138498 407086
rect 139301 407083 139367 407086
rect 150934 407084 150940 407148
rect 151004 407146 151010 407148
rect 151353 407146 151419 407149
rect 151004 407144 151419 407146
rect 151004 407088 151358 407144
rect 151414 407088 151419 407144
rect 151004 407086 151419 407088
rect 151004 407084 151010 407086
rect 151353 407083 151419 407086
rect 208710 407084 208716 407148
rect 208780 407146 208786 407148
rect 209497 407146 209563 407149
rect 211061 407148 211127 407149
rect 211061 407146 211108 407148
rect 208780 407144 209563 407146
rect 208780 407088 209502 407144
rect 209558 407088 209563 407144
rect 208780 407086 209563 407088
rect 211016 407144 211108 407146
rect 211016 407088 211066 407144
rect 211016 407086 211108 407088
rect 208780 407084 208786 407086
rect 209497 407083 209563 407086
rect 211061 407084 211108 407086
rect 211172 407084 211178 407148
rect 218462 407084 218468 407148
rect 218532 407146 218538 407148
rect 218973 407146 219039 407149
rect 218532 407144 219039 407146
rect 218532 407088 218978 407144
rect 219034 407088 219039 407144
rect 218532 407086 219039 407088
rect 218532 407084 218538 407086
rect 211061 407083 211127 407084
rect 218973 407083 219039 407086
rect 231158 407084 231164 407148
rect 231228 407146 231234 407148
rect 231761 407146 231827 407149
rect 231228 407144 231827 407146
rect 231228 407088 231766 407144
rect 231822 407088 231827 407144
rect 231228 407086 231827 407088
rect 231228 407084 231234 407086
rect 231761 407083 231827 407086
rect 233550 407084 233556 407148
rect 233620 407146 233626 407148
rect 234521 407146 234587 407149
rect 233620 407144 234587 407146
rect 233620 407088 234526 407144
rect 234582 407088 234587 407144
rect 233620 407086 234587 407088
rect 233620 407084 233626 407086
rect 234521 407083 234587 407086
rect 236126 407084 236132 407148
rect 236196 407146 236202 407148
rect 237281 407146 237347 407149
rect 236196 407144 237347 407146
rect 236196 407088 237286 407144
rect 237342 407088 237347 407144
rect 236196 407086 237347 407088
rect 236196 407084 236202 407086
rect 237281 407083 237347 407086
rect 240910 407084 240916 407148
rect 240980 407146 240986 407148
rect 241421 407146 241487 407149
rect 240980 407144 241487 407146
rect 240980 407088 241426 407144
rect 241482 407088 241487 407144
rect 240980 407086 241487 407088
rect 240980 407084 240986 407086
rect 241421 407083 241487 407086
rect 246062 407084 246068 407148
rect 246132 407146 246138 407148
rect 246941 407146 247007 407149
rect 246132 407144 247007 407146
rect 246132 407088 246946 407144
rect 247002 407088 247007 407144
rect 246132 407086 247007 407088
rect 246132 407084 246138 407086
rect 246941 407083 247007 407086
rect 248638 407084 248644 407148
rect 248708 407146 248714 407148
rect 249701 407146 249767 407149
rect 248708 407144 249767 407146
rect 248708 407088 249706 407144
rect 249762 407088 249767 407144
rect 248708 407086 249767 407088
rect 248708 407084 248714 407086
rect 249701 407083 249767 407086
rect 255998 407084 256004 407148
rect 256068 407146 256074 407148
rect 256601 407146 256667 407149
rect 256068 407144 256667 407146
rect 256068 407088 256606 407144
rect 256662 407088 256667 407144
rect 256068 407086 256667 407088
rect 256068 407084 256074 407086
rect 256601 407083 256667 407086
rect 261150 407084 261156 407148
rect 261220 407146 261226 407148
rect 262121 407146 262187 407149
rect 261220 407144 262187 407146
rect 261220 407088 262126 407144
rect 262182 407088 262187 407144
rect 261220 407086 262187 407088
rect 261220 407084 261226 407086
rect 262121 407083 262187 407086
rect 276054 407084 276060 407148
rect 276124 407146 276130 407148
rect 276841 407146 276907 407149
rect 276124 407144 276907 407146
rect 276124 407088 276846 407144
rect 276902 407088 276907 407144
rect 276124 407086 276907 407088
rect 276124 407084 276130 407086
rect 276841 407083 276907 407086
rect 283414 407084 283420 407148
rect 283484 407146 283490 407148
rect 284201 407146 284267 407149
rect 283484 407144 284267 407146
rect 283484 407088 284206 407144
rect 284262 407088 284267 407144
rect 283484 407086 284267 407088
rect 283484 407084 283490 407086
rect 284201 407083 284267 407086
rect 298502 407084 298508 407148
rect 298572 407146 298578 407148
rect 299381 407146 299447 407149
rect 298572 407144 299447 407146
rect 298572 407088 299386 407144
rect 299442 407088 299447 407144
rect 298572 407086 299447 407088
rect 298572 407084 298578 407086
rect 299381 407083 299447 407086
rect 299790 407084 299796 407148
rect 299860 407146 299866 407148
rect 300761 407146 300827 407149
rect 299860 407144 300827 407146
rect 299860 407088 300766 407144
rect 300822 407088 300827 407144
rect 299860 407086 300827 407088
rect 299860 407084 299866 407086
rect 300761 407083 300827 407086
rect 310830 407084 310836 407148
rect 310900 407146 310906 407148
rect 317413 407146 317479 407149
rect 310900 407144 317479 407146
rect 310900 407088 317418 407144
rect 317474 407088 317479 407144
rect 310900 407086 317479 407088
rect 310900 407084 310906 407086
rect 317413 407083 317479 407086
rect 86217 406604 86283 406605
rect 88609 406604 88675 406605
rect 95969 406604 96035 406605
rect 238569 406604 238635 406605
rect 243721 406604 243787 406605
rect 281073 406604 281139 406605
rect 78438 406540 78444 406604
rect 78508 406602 78514 406604
rect 78508 406542 84210 406602
rect 78508 406540 78514 406542
rect 81065 406468 81131 406469
rect 83641 406468 83707 406469
rect 81014 406404 81020 406468
rect 81084 406466 81131 406468
rect 81084 406464 81176 406466
rect 81126 406408 81176 406464
rect 81084 406406 81176 406408
rect 81084 406404 81131 406406
rect 83590 406404 83596 406468
rect 83660 406466 83707 406468
rect 84150 406466 84210 406542
rect 86166 406540 86172 406604
rect 86236 406602 86283 406604
rect 86236 406600 86328 406602
rect 86278 406544 86328 406600
rect 86236 406542 86328 406544
rect 86236 406540 86283 406542
rect 88558 406540 88564 406604
rect 88628 406602 88675 406604
rect 88628 406600 88720 406602
rect 88670 406544 88720 406600
rect 88628 406542 88720 406544
rect 88628 406540 88675 406542
rect 95918 406540 95924 406604
rect 95988 406602 96035 406604
rect 95988 406600 96080 406602
rect 96030 406544 96080 406600
rect 95988 406542 96080 406544
rect 95988 406540 96035 406542
rect 238518 406540 238524 406604
rect 238588 406602 238635 406604
rect 238588 406600 238680 406602
rect 238630 406544 238680 406600
rect 238588 406542 238680 406544
rect 238588 406540 238635 406542
rect 243670 406540 243676 406604
rect 243740 406602 243787 406604
rect 243740 406600 243832 406602
rect 243782 406544 243832 406600
rect 243740 406542 243832 406544
rect 243740 406540 243787 406542
rect 281022 406540 281028 406604
rect 281092 406602 281139 406604
rect 281092 406600 281184 406602
rect 281134 406544 281184 406600
rect 281092 406542 281184 406544
rect 281092 406540 281139 406542
rect 86217 406539 86283 406540
rect 88609 406539 88675 406540
rect 95969 406539 96035 406540
rect 238569 406539 238635 406540
rect 243721 406539 243787 406540
rect 281073 406539 281139 406540
rect 325233 406466 325299 406469
rect 83660 406464 83752 406466
rect 83702 406408 83752 406464
rect 83660 406406 83752 406408
rect 84150 406464 325299 406466
rect 84150 406408 325238 406464
rect 325294 406408 325299 406464
rect 84150 406406 325299 406408
rect 83660 406404 83707 406406
rect 81065 406403 81131 406404
rect 83641 406403 83707 406404
rect 325233 406403 325299 406406
rect 321093 406330 321159 406333
rect 74490 406328 321159 406330
rect 74490 406272 321098 406328
rect 321154 406272 321159 406328
rect 74490 406270 321159 406272
rect 48681 406196 48747 406197
rect 53465 406196 53531 406197
rect 61101 406196 61167 406197
rect 48681 406194 48702 406196
rect 48610 406192 48702 406194
rect 48610 406136 48686 406192
rect 48610 406134 48702 406136
rect 48681 406132 48702 406134
rect 48766 406132 48772 406196
rect 53456 406132 53462 406196
rect 53526 406194 53532 406196
rect 53526 406134 53618 406194
rect 53526 406132 53532 406134
rect 61072 406132 61078 406196
rect 61142 406194 61167 406196
rect 61142 406192 61234 406194
rect 61162 406136 61234 406192
rect 61142 406134 61234 406136
rect 61142 406132 61167 406134
rect 73584 406132 73590 406196
rect 73654 406194 73660 406196
rect 74490 406194 74550 406270
rect 321093 406267 321159 406270
rect 73654 406134 74550 406194
rect 73654 406132 73660 406134
rect 76168 406132 76174 406196
rect 76238 406194 76244 406196
rect 330661 406194 330727 406197
rect 76238 406192 330727 406194
rect 76238 406136 330666 406192
rect 330722 406136 330727 406192
rect 76238 406134 330727 406136
rect 76238 406132 76244 406134
rect 48681 406131 48747 406132
rect 53465 406131 53531 406132
rect 61101 406131 61167 406132
rect 330661 406131 330727 406134
rect 3601 406058 3667 406061
rect 316861 406058 316927 406061
rect 3601 406056 316927 406058
rect 3601 406000 3606 406056
rect 3662 406000 316866 406056
rect 316922 406000 316927 406056
rect 3601 405998 316927 406000
rect 3601 405995 3667 405998
rect 316861 405995 316927 405998
rect 3417 405922 3483 405925
rect 318149 405922 318215 405925
rect 3417 405920 318215 405922
rect 3417 405864 3422 405920
rect 3478 405864 318154 405920
rect 318210 405864 318215 405920
rect 3417 405862 318215 405864
rect 3417 405859 3483 405862
rect 318149 405859 318215 405862
rect 583520 404820 584960 405060
rect 159357 401706 159423 401709
rect 320081 401706 320147 401709
rect 157198 401704 159423 401706
rect 157198 401648 159362 401704
rect 159418 401648 159423 401704
rect 157198 401646 159423 401648
rect 157198 401620 157258 401646
rect 159357 401643 159423 401646
rect 317094 401704 320147 401706
rect 317094 401648 320086 401704
rect 320142 401648 320147 401704
rect 317094 401646 320147 401648
rect 317094 401620 317154 401646
rect 320081 401643 320147 401646
rect 156588 401560 157258 401620
rect 316572 401560 317154 401620
rect 337653 397626 337719 397629
rect 337653 397624 340124 397626
rect -960 397490 480 397580
rect 337653 397568 337658 397624
rect 337714 397568 340124 397624
rect 337653 397566 340124 397568
rect 337653 397563 337719 397566
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 337653 396946 337719 396949
rect 337653 396944 340124 396946
rect 337653 396888 337658 396944
rect 337714 396888 340124 396944
rect 337653 396886 340124 396888
rect 337653 396883 337719 396886
rect 335997 396266 336063 396269
rect 335997 396264 340124 396266
rect 335997 396208 336002 396264
rect 336058 396208 340124 396264
rect 335997 396206 340124 396208
rect 335997 396203 336063 396206
rect 337745 395722 337811 395725
rect 337745 395720 340124 395722
rect 337745 395664 337750 395720
rect 337806 395664 340124 395720
rect 337745 395662 340124 395664
rect 337745 395659 337811 395662
rect 482921 395586 482987 395589
rect 479964 395584 482987 395586
rect 479964 395528 482926 395584
rect 482982 395528 482987 395584
rect 479964 395526 482987 395528
rect 482921 395523 482987 395526
rect 337653 395042 337719 395045
rect 337653 395040 340124 395042
rect 337653 394984 337658 395040
rect 337714 394984 340124 395040
rect 337653 394982 340124 394984
rect 337653 394979 337719 394982
rect 337745 394362 337811 394365
rect 337745 394360 340124 394362
rect 337745 394304 337750 394360
rect 337806 394304 340124 394360
rect 337745 394302 340124 394304
rect 337745 394299 337811 394302
rect 337653 393682 337719 393685
rect 337653 393680 340124 393682
rect 337653 393624 337658 393680
rect 337714 393624 340124 393680
rect 337653 393622 340124 393624
rect 337653 393619 337719 393622
rect 337745 393138 337811 393141
rect 337745 393136 340124 393138
rect 337745 393080 337750 393136
rect 337806 393080 340124 393136
rect 337745 393078 340124 393080
rect 337745 393075 337811 393078
rect 337653 392458 337719 392461
rect 337653 392456 340124 392458
rect 337653 392400 337658 392456
rect 337714 392400 340124 392456
rect 337653 392398 340124 392400
rect 337653 392395 337719 392398
rect 337653 391778 337719 391781
rect 337653 391776 340124 391778
rect 337653 391720 337658 391776
rect 337714 391720 340124 391776
rect 337653 391718 340124 391720
rect 337653 391715 337719 391718
rect 583520 391628 584960 391868
rect 337745 391234 337811 391237
rect 337745 391232 340124 391234
rect 337745 391176 337750 391232
rect 337806 391176 340124 391232
rect 337745 391174 340124 391176
rect 337745 391171 337811 391174
rect 482921 390962 482987 390965
rect 479964 390960 482987 390962
rect 479964 390904 482926 390960
rect 482982 390904 482987 390960
rect 479964 390902 482987 390904
rect 482921 390899 482987 390902
rect 337653 390554 337719 390557
rect 337653 390552 340124 390554
rect 337653 390496 337658 390552
rect 337714 390496 340124 390552
rect 337653 390494 340124 390496
rect 337653 390491 337719 390494
rect 337745 389874 337811 389877
rect 337745 389872 340124 389874
rect 337745 389816 337750 389872
rect 337806 389816 340124 389872
rect 337745 389814 340124 389816
rect 337745 389811 337811 389814
rect 337653 389194 337719 389197
rect 337653 389192 340124 389194
rect 337653 389136 337658 389192
rect 337714 389136 340124 389192
rect 337653 389134 340124 389136
rect 337653 389131 337719 389134
rect 337745 388650 337811 388653
rect 337745 388648 340124 388650
rect 337745 388592 337750 388648
rect 337806 388592 340124 388648
rect 337745 388590 340124 388592
rect 337745 388587 337811 388590
rect 337837 387970 337903 387973
rect 337837 387968 340124 387970
rect 337837 387912 337842 387968
rect 337898 387912 340124 387968
rect 337837 387910 340124 387912
rect 337837 387907 337903 387910
rect 337653 387290 337719 387293
rect 337653 387288 340124 387290
rect 337653 387232 337658 387288
rect 337714 387232 340124 387288
rect 337653 387230 340124 387232
rect 337653 387227 337719 387230
rect 337745 386746 337811 386749
rect 337745 386744 340124 386746
rect 337745 386688 337750 386744
rect 337806 386688 340124 386744
rect 337745 386686 340124 386688
rect 337745 386683 337811 386686
rect 482921 386338 482987 386341
rect 479964 386336 482987 386338
rect 479964 386280 482926 386336
rect 482982 386280 482987 386336
rect 479964 386278 482987 386280
rect 482921 386275 482987 386278
rect 337653 386066 337719 386069
rect 337653 386064 340124 386066
rect 337653 386008 337658 386064
rect 337714 386008 340124 386064
rect 337653 386006 340124 386008
rect 337653 386003 337719 386006
rect 337745 385386 337811 385389
rect 337745 385384 340124 385386
rect 337745 385328 337750 385384
rect 337806 385328 340124 385384
rect 337745 385326 340124 385328
rect 337745 385323 337811 385326
rect 337653 384706 337719 384709
rect 337653 384704 340124 384706
rect 337653 384648 337658 384704
rect 337714 384648 340124 384704
rect 337653 384646 340124 384648
rect 337653 384643 337719 384646
rect -960 384284 480 384524
rect 337745 384162 337811 384165
rect 337745 384160 340124 384162
rect 337745 384104 337750 384160
rect 337806 384104 340124 384160
rect 337745 384102 340124 384104
rect 337745 384099 337811 384102
rect 337653 383482 337719 383485
rect 337653 383480 340124 383482
rect 337653 383424 337658 383480
rect 337714 383424 340124 383480
rect 337653 383422 340124 383424
rect 337653 383419 337719 383422
rect 337745 382802 337811 382805
rect 337745 382800 340124 382802
rect 337745 382744 337750 382800
rect 337806 382744 340124 382800
rect 337745 382742 340124 382744
rect 337745 382739 337811 382742
rect 337653 382122 337719 382125
rect 337653 382120 340124 382122
rect 337653 382064 337658 382120
rect 337714 382064 340124 382120
rect 337653 382062 340124 382064
rect 337653 382059 337719 382062
rect 336917 381578 336983 381581
rect 482001 381578 482067 381581
rect 336917 381576 340124 381578
rect 336917 381520 336922 381576
rect 336978 381520 340124 381576
rect 336917 381518 340124 381520
rect 479964 381576 482067 381578
rect 479964 381520 482006 381576
rect 482062 381520 482067 381576
rect 479964 381518 482067 381520
rect 336917 381515 336983 381518
rect 482001 381515 482067 381518
rect 336089 380898 336155 380901
rect 336089 380896 340124 380898
rect 336089 380840 336094 380896
rect 336150 380840 340124 380896
rect 336089 380838 340124 380840
rect 336089 380835 336155 380838
rect 337745 380218 337811 380221
rect 337745 380216 340124 380218
rect 337745 380160 337750 380216
rect 337806 380160 340124 380216
rect 337745 380158 340124 380160
rect 337745 380155 337811 380158
rect 336917 379674 336983 379677
rect 336917 379672 340124 379674
rect 336917 379616 336922 379672
rect 336978 379616 340124 379672
rect 336917 379614 340124 379616
rect 336917 379611 336983 379614
rect 337653 378994 337719 378997
rect 337653 378992 340124 378994
rect 337653 378936 337658 378992
rect 337714 378936 340124 378992
rect 337653 378934 340124 378936
rect 337653 378931 337719 378934
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 337745 378314 337811 378317
rect 337745 378312 340124 378314
rect 337745 378256 337750 378312
rect 337806 378256 340124 378312
rect 583520 378300 584960 378390
rect 337745 378254 340124 378256
rect 337745 378251 337811 378254
rect 337285 377634 337351 377637
rect 337285 377632 340124 377634
rect 337285 377576 337290 377632
rect 337346 377576 340124 377632
rect 337285 377574 340124 377576
rect 337285 377571 337351 377574
rect 337745 377090 337811 377093
rect 337745 377088 340124 377090
rect 337745 377032 337750 377088
rect 337806 377032 340124 377088
rect 337745 377030 340124 377032
rect 337745 377027 337811 377030
rect 482277 376954 482343 376957
rect 479964 376952 482343 376954
rect 479964 376896 482282 376952
rect 482338 376896 482343 376952
rect 479964 376894 482343 376896
rect 482277 376891 482343 376894
rect 337101 376410 337167 376413
rect 337101 376408 340124 376410
rect 337101 376352 337106 376408
rect 337162 376352 340124 376408
rect 337101 376350 340124 376352
rect 337101 376347 337167 376350
rect 337653 375730 337719 375733
rect 337653 375728 340124 375730
rect 337653 375672 337658 375728
rect 337714 375672 340124 375728
rect 337653 375670 340124 375672
rect 337653 375667 337719 375670
rect 337745 375186 337811 375189
rect 337745 375184 340124 375186
rect 337745 375128 337750 375184
rect 337806 375128 340124 375184
rect 337745 375126 340124 375128
rect 337745 375123 337811 375126
rect 337653 374506 337719 374509
rect 337653 374504 340124 374506
rect 337653 374448 337658 374504
rect 337714 374448 340124 374504
rect 337653 374446 340124 374448
rect 337653 374443 337719 374446
rect 337745 373826 337811 373829
rect 337745 373824 340124 373826
rect 337745 373768 337750 373824
rect 337806 373768 340124 373824
rect 337745 373766 340124 373768
rect 337745 373763 337811 373766
rect 337653 373146 337719 373149
rect 337653 373144 340124 373146
rect 337653 373088 337658 373144
rect 337714 373088 340124 373144
rect 337653 373086 340124 373088
rect 337653 373083 337719 373086
rect 336917 372602 336983 372605
rect 336917 372600 340124 372602
rect 336917 372544 336922 372600
rect 336978 372544 340124 372600
rect 336917 372542 340124 372544
rect 336917 372539 336983 372542
rect 482921 372330 482987 372333
rect 479964 372328 482987 372330
rect 479964 372272 482926 372328
rect 482982 372272 482987 372328
rect 479964 372270 482987 372272
rect 482921 372267 482987 372270
rect 337561 371922 337627 371925
rect 337561 371920 340124 371922
rect 337561 371864 337566 371920
rect 337622 371864 340124 371920
rect 337561 371862 340124 371864
rect 337561 371859 337627 371862
rect -960 371228 480 371468
rect 336457 371242 336523 371245
rect 336457 371240 340124 371242
rect 336457 371184 336462 371240
rect 336518 371184 340124 371240
rect 336457 371182 340124 371184
rect 336457 371179 336523 371182
rect 337653 370698 337719 370701
rect 337653 370696 340124 370698
rect 337653 370640 337658 370696
rect 337714 370640 340124 370696
rect 337653 370638 340124 370640
rect 337653 370635 337719 370638
rect 337653 370018 337719 370021
rect 337653 370016 340124 370018
rect 337653 369960 337658 370016
rect 337714 369960 340124 370016
rect 337653 369958 340124 369960
rect 337653 369955 337719 369958
rect 337285 369338 337351 369341
rect 337285 369336 340124 369338
rect 337285 369280 337290 369336
rect 337346 369280 340124 369336
rect 337285 369278 340124 369280
rect 337285 369275 337351 369278
rect 337653 368658 337719 368661
rect 337653 368656 340124 368658
rect 337653 368600 337658 368656
rect 337714 368600 340124 368656
rect 337653 368598 340124 368600
rect 337653 368595 337719 368598
rect 337745 368114 337811 368117
rect 337745 368112 340124 368114
rect 337745 368056 337750 368112
rect 337806 368056 340124 368112
rect 337745 368054 340124 368056
rect 337745 368051 337811 368054
rect 482369 367570 482435 367573
rect 479964 367568 482435 367570
rect 479964 367512 482374 367568
rect 482430 367512 482435 367568
rect 479964 367510 482435 367512
rect 482369 367507 482435 367510
rect 337745 367434 337811 367437
rect 337745 367432 340124 367434
rect 337745 367376 337750 367432
rect 337806 367376 340124 367432
rect 337745 367374 340124 367376
rect 337745 367371 337811 367374
rect 336549 366754 336615 366757
rect 336549 366752 340124 366754
rect 336549 366696 336554 366752
rect 336610 366696 340124 366752
rect 336549 366694 340124 366696
rect 336549 366691 336615 366694
rect 337285 366074 337351 366077
rect 337285 366072 340124 366074
rect 337285 366016 337290 366072
rect 337346 366016 340124 366072
rect 337285 366014 340124 366016
rect 337285 366011 337351 366014
rect 337653 365530 337719 365533
rect 337653 365528 340124 365530
rect 337653 365472 337658 365528
rect 337714 365472 340124 365528
rect 337653 365470 340124 365472
rect 337653 365467 337719 365470
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 337745 364850 337811 364853
rect 337745 364848 340124 364850
rect 337745 364792 337750 364848
rect 337806 364792 340124 364848
rect 337745 364790 340124 364792
rect 337745 364787 337811 364790
rect 337653 364170 337719 364173
rect 337653 364168 340124 364170
rect 337653 364112 337658 364168
rect 337714 364112 340124 364168
rect 337653 364110 340124 364112
rect 337653 364107 337719 364110
rect 337745 363626 337811 363629
rect 337745 363624 340124 363626
rect 337745 363568 337750 363624
rect 337806 363568 340124 363624
rect 337745 363566 340124 363568
rect 337745 363563 337811 363566
rect 337653 362946 337719 362949
rect 482461 362946 482527 362949
rect 337653 362944 340124 362946
rect 337653 362888 337658 362944
rect 337714 362888 340124 362944
rect 337653 362886 340124 362888
rect 479964 362944 482527 362946
rect 479964 362888 482466 362944
rect 482522 362888 482527 362944
rect 479964 362886 482527 362888
rect 337653 362883 337719 362886
rect 482461 362883 482527 362886
rect 337101 362266 337167 362269
rect 337101 362264 340124 362266
rect 337101 362208 337106 362264
rect 337162 362208 340124 362264
rect 337101 362206 340124 362208
rect 337101 362203 337167 362206
rect 337561 361586 337627 361589
rect 337561 361584 340124 361586
rect 337561 361528 337566 361584
rect 337622 361528 340124 361584
rect 337561 361526 340124 361528
rect 337561 361523 337627 361526
rect 337653 361042 337719 361045
rect 337653 361040 340124 361042
rect 337653 360984 337658 361040
rect 337714 360984 340124 361040
rect 337653 360982 340124 360984
rect 337653 360979 337719 360982
rect 336917 360362 336983 360365
rect 336917 360360 340124 360362
rect 336917 360304 336922 360360
rect 336978 360304 340124 360360
rect 336917 360302 340124 360304
rect 336917 360299 336983 360302
rect 337653 359682 337719 359685
rect 337653 359680 340124 359682
rect 337653 359624 337658 359680
rect 337714 359624 340124 359680
rect 337653 359622 340124 359624
rect 337653 359619 337719 359622
rect 17125 359274 17191 359277
rect 19382 359274 20056 359324
rect 17125 359272 20056 359274
rect 17125 359216 17130 359272
rect 17186 359264 20056 359272
rect 177205 359274 177271 359277
rect 179462 359274 180032 359324
rect 177205 359272 180032 359274
rect 17186 359216 19442 359264
rect 17125 359214 19442 359216
rect 177205 359216 177210 359272
rect 177266 359264 180032 359272
rect 177266 359216 179522 359264
rect 177205 359214 179522 359216
rect 17125 359211 17191 359214
rect 177205 359211 177271 359214
rect 337469 359138 337535 359141
rect 337469 359136 340124 359138
rect 337469 359080 337474 359136
rect 337530 359080 340124 359136
rect 337469 359078 340124 359080
rect 337469 359075 337535 359078
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 337745 358458 337811 358461
rect 337745 358456 340124 358458
rect 337745 358400 337750 358456
rect 337806 358400 340124 358456
rect 337745 358398 340124 358400
rect 337745 358395 337811 358398
rect 17217 358322 17283 358325
rect 19382 358322 20056 358372
rect 17217 358320 20056 358322
rect 17217 358264 17222 358320
rect 17278 358312 20056 358320
rect 177389 358322 177455 358325
rect 179462 358322 180032 358372
rect 482553 358322 482619 358325
rect 177389 358320 180032 358322
rect 17278 358264 19442 358312
rect 17217 358262 19442 358264
rect 177389 358264 177394 358320
rect 177450 358312 180032 358320
rect 479964 358320 482619 358322
rect 177450 358264 179522 358312
rect 177389 358262 179522 358264
rect 479964 358264 482558 358320
rect 482614 358264 482619 358320
rect 479964 358262 482619 358264
rect 17217 358259 17283 358262
rect 177389 358259 177455 358262
rect 482553 358259 482619 358262
rect 336917 357778 336983 357781
rect 336917 357776 340124 357778
rect 336917 357720 336922 357776
rect 336978 357720 340124 357776
rect 336917 357718 340124 357720
rect 336917 357715 336983 357718
rect 336089 357098 336155 357101
rect 336089 357096 340124 357098
rect 336089 357040 336094 357096
rect 336150 357040 340124 357096
rect 336089 357038 340124 357040
rect 336089 357035 336155 357038
rect 337653 356554 337719 356557
rect 337653 356552 340124 356554
rect 337653 356496 337658 356552
rect 337714 356496 340124 356552
rect 337653 356494 340124 356496
rect 337653 356491 337719 356494
rect 17769 356146 17835 356149
rect 19382 356146 20056 356196
rect 17769 356144 20056 356146
rect 17769 356088 17774 356144
rect 17830 356136 20056 356144
rect 177849 356146 177915 356149
rect 179462 356146 180032 356196
rect 177849 356144 180032 356146
rect 17830 356088 19442 356136
rect 17769 356086 19442 356088
rect 177849 356088 177854 356144
rect 177910 356136 180032 356144
rect 177910 356088 179522 356136
rect 177849 356086 179522 356088
rect 17769 356083 17835 356086
rect 177849 356083 177915 356086
rect 337653 355874 337719 355877
rect 337653 355872 340124 355874
rect 337653 355816 337658 355872
rect 337714 355816 340124 355872
rect 337653 355814 340124 355816
rect 337653 355811 337719 355814
rect 17677 355194 17743 355197
rect 19382 355194 20056 355244
rect 17677 355192 20056 355194
rect 17677 355136 17682 355192
rect 17738 355184 20056 355192
rect 177757 355194 177823 355197
rect 179462 355194 180032 355244
rect 177757 355192 180032 355194
rect 17738 355136 19442 355184
rect 17677 355134 19442 355136
rect 177757 355136 177762 355192
rect 177818 355184 180032 355192
rect 336365 355194 336431 355197
rect 336365 355192 340124 355194
rect 177818 355136 179522 355184
rect 177757 355134 179522 355136
rect 336365 355136 336370 355192
rect 336426 355136 340124 355192
rect 336365 355134 340124 355136
rect 17677 355131 17743 355134
rect 177757 355131 177823 355134
rect 336365 355131 336431 355134
rect 337745 354650 337811 354653
rect 337745 354648 340124 354650
rect 337745 354592 337750 354648
rect 337806 354592 340124 354648
rect 337745 354590 340124 354592
rect 337745 354587 337811 354590
rect 337561 353970 337627 353973
rect 337561 353968 340124 353970
rect 337561 353912 337566 353968
rect 337622 353912 340124 353968
rect 337561 353910 340124 353912
rect 337561 353907 337627 353910
rect 482645 353698 482711 353701
rect 479964 353696 482711 353698
rect 479964 353640 482650 353696
rect 482706 353640 482711 353696
rect 479964 353638 482711 353640
rect 482645 353635 482711 353638
rect 17493 353426 17559 353429
rect 19382 353426 20056 353476
rect 17493 353424 20056 353426
rect 17493 353368 17498 353424
rect 17554 353416 20056 353424
rect 177665 353426 177731 353429
rect 179462 353426 180032 353476
rect 177665 353424 180032 353426
rect 17554 353368 19442 353416
rect 17493 353366 19442 353368
rect 177665 353368 177670 353424
rect 177726 353416 180032 353424
rect 177726 353368 179522 353416
rect 177665 353366 179522 353368
rect 17493 353363 17559 353366
rect 177665 353363 177731 353366
rect 336917 353290 336983 353293
rect 336917 353288 340124 353290
rect 336917 353232 336922 353288
rect 336978 353232 340124 353288
rect 336917 353230 340124 353232
rect 336917 353227 336983 353230
rect 337653 352610 337719 352613
rect 337653 352608 340124 352610
rect 337653 352552 337658 352608
rect 337714 352552 340124 352608
rect 337653 352550 340124 352552
rect 337653 352547 337719 352550
rect 17401 352338 17467 352341
rect 19382 352338 20056 352388
rect 17401 352336 20056 352338
rect 17401 352280 17406 352336
rect 17462 352328 20056 352336
rect 177573 352338 177639 352341
rect 179462 352338 180032 352388
rect 177573 352336 180032 352338
rect 17462 352280 19442 352328
rect 17401 352278 19442 352280
rect 177573 352280 177578 352336
rect 177634 352328 180032 352336
rect 177634 352280 179522 352328
rect 177573 352278 179522 352280
rect 17401 352275 17467 352278
rect 177573 352275 177639 352278
rect 337285 352066 337351 352069
rect 337285 352064 340124 352066
rect 337285 352008 337290 352064
rect 337346 352008 340124 352064
rect 337285 352006 340124 352008
rect 337285 352003 337351 352006
rect 583520 351780 584960 352020
rect 337653 351386 337719 351389
rect 337653 351384 340124 351386
rect 337653 351328 337658 351384
rect 337714 351328 340124 351384
rect 337653 351326 340124 351328
rect 337653 351323 337719 351326
rect 337653 350706 337719 350709
rect 337653 350704 340124 350706
rect 337653 350648 337658 350704
rect 337714 350648 340124 350704
rect 337653 350646 340124 350648
rect 337653 350643 337719 350646
rect 17585 350570 17651 350573
rect 19382 350570 20056 350620
rect 17585 350568 20056 350570
rect 17585 350512 17590 350568
rect 17646 350560 20056 350568
rect 177481 350570 177547 350573
rect 179462 350570 180032 350620
rect 177481 350568 180032 350570
rect 17646 350512 19442 350560
rect 17585 350510 19442 350512
rect 177481 350512 177486 350568
rect 177542 350560 180032 350568
rect 177542 350512 179522 350560
rect 177481 350510 179522 350512
rect 17585 350507 17651 350510
rect 177481 350507 177547 350510
rect 337745 350026 337811 350029
rect 337745 350024 340124 350026
rect 337745 349968 337750 350024
rect 337806 349968 340124 350024
rect 337745 349966 340124 349968
rect 337745 349963 337811 349966
rect 337653 349482 337719 349485
rect 337653 349480 340124 349482
rect 337653 349424 337658 349480
rect 337714 349424 340124 349480
rect 337653 349422 340124 349424
rect 337653 349419 337719 349422
rect 482737 348938 482803 348941
rect 479964 348936 482803 348938
rect 479964 348880 482742 348936
rect 482798 348880 482803 348936
rect 479964 348878 482803 348880
rect 482737 348875 482803 348878
rect 337745 348802 337811 348805
rect 337745 348800 340124 348802
rect 337745 348744 337750 348800
rect 337806 348744 340124 348800
rect 337745 348742 340124 348744
rect 337745 348739 337811 348742
rect 336365 348122 336431 348125
rect 336365 348120 340124 348122
rect 336365 348064 336370 348120
rect 336426 348064 340124 348120
rect 336365 348062 340124 348064
rect 336365 348059 336431 348062
rect 337653 347578 337719 347581
rect 337653 347576 340124 347578
rect 337653 347520 337658 347576
rect 337714 347520 340124 347576
rect 337653 347518 340124 347520
rect 337653 347515 337719 347518
rect 337469 346898 337535 346901
rect 337469 346896 340124 346898
rect 337469 346840 337474 346896
rect 337530 346840 340124 346896
rect 337469 346838 340124 346840
rect 337469 346835 337535 346838
rect 337653 346218 337719 346221
rect 337653 346216 340124 346218
rect 337653 346160 337658 346216
rect 337714 346160 340124 346216
rect 337653 346158 340124 346160
rect 337653 346155 337719 346158
rect 337653 345538 337719 345541
rect 337653 345536 340124 345538
rect -960 345402 480 345492
rect 337653 345480 337658 345536
rect 337714 345480 340124 345536
rect 337653 345478 340124 345480
rect 337653 345475 337719 345478
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 337745 344994 337811 344997
rect 337745 344992 340124 344994
rect 337745 344936 337750 344992
rect 337806 344936 340124 344992
rect 337745 344934 340124 344936
rect 337745 344931 337811 344934
rect 337653 344314 337719 344317
rect 482829 344314 482895 344317
rect 337653 344312 340124 344314
rect 337653 344256 337658 344312
rect 337714 344256 340124 344312
rect 337653 344254 340124 344256
rect 479964 344312 482895 344314
rect 479964 344256 482834 344312
rect 482890 344256 482895 344312
rect 479964 344254 482895 344256
rect 337653 344251 337719 344254
rect 482829 344251 482895 344254
rect 337745 343634 337811 343637
rect 337745 343632 340124 343634
rect 337745 343576 337750 343632
rect 337806 343576 340124 343632
rect 337745 343574 340124 343576
rect 337745 343571 337811 343574
rect 337653 343090 337719 343093
rect 337653 343088 340124 343090
rect 337653 343032 337658 343088
rect 337714 343032 340124 343088
rect 337653 343030 340124 343032
rect 337653 343027 337719 343030
rect 337561 342410 337627 342413
rect 337561 342408 340124 342410
rect 337561 342352 337566 342408
rect 337622 342352 340124 342408
rect 337561 342350 340124 342352
rect 337561 342347 337627 342350
rect 156588 341730 157258 341780
rect 159081 341730 159147 341733
rect 156588 341728 159147 341730
rect 156588 341720 159086 341728
rect 157198 341672 159086 341720
rect 159142 341672 159147 341728
rect 316572 341730 317154 341780
rect 319529 341730 319595 341733
rect 316572 341728 319595 341730
rect 316572 341720 319534 341728
rect 157198 341670 159147 341672
rect 317094 341672 319534 341720
rect 319590 341672 319595 341728
rect 317094 341670 319595 341672
rect 159081 341667 159147 341670
rect 319529 341667 319595 341670
rect 336273 341730 336339 341733
rect 336273 341728 340124 341730
rect 336273 341672 336278 341728
rect 336334 341672 340124 341728
rect 336273 341670 340124 341672
rect 336273 341667 336339 341670
rect 336917 341050 336983 341053
rect 336917 341048 340124 341050
rect 336917 340992 336922 341048
rect 336978 340992 340124 341048
rect 336917 340990 340124 340992
rect 336917 340987 336983 340990
rect 337285 340506 337351 340509
rect 337285 340504 340124 340506
rect 337285 340448 337290 340504
rect 337346 340448 340124 340504
rect 337285 340446 340124 340448
rect 337285 340443 337351 340446
rect 156588 340098 157258 340148
rect 158713 340098 158779 340101
rect 156588 340096 158779 340098
rect 156588 340088 158718 340096
rect 157198 340040 158718 340088
rect 158774 340040 158779 340096
rect 316572 340098 317154 340148
rect 319621 340098 319687 340101
rect 316572 340096 319687 340098
rect 316572 340088 319626 340096
rect 157198 340038 158779 340040
rect 317094 340040 319626 340088
rect 319682 340040 319687 340096
rect 317094 340038 319687 340040
rect 158713 340035 158779 340038
rect 319621 340035 319687 340038
rect 336181 339826 336247 339829
rect 336181 339824 340124 339826
rect 336181 339768 336186 339824
rect 336242 339768 340124 339824
rect 336181 339766 340124 339768
rect 336181 339763 336247 339766
rect 482277 339690 482343 339693
rect 479964 339688 482343 339690
rect 479964 339632 482282 339688
rect 482338 339632 482343 339688
rect 479964 339630 482343 339632
rect 482277 339627 482343 339630
rect 337285 339146 337351 339149
rect 337285 339144 340124 339146
rect 337285 339088 337290 339144
rect 337346 339088 340124 339144
rect 337285 339086 340124 339088
rect 337285 339083 337351 339086
rect 156588 338738 157258 338788
rect 158805 338738 158871 338741
rect 156588 338736 158871 338738
rect 156588 338728 158810 338736
rect 157198 338680 158810 338728
rect 158866 338680 158871 338736
rect 316572 338738 317154 338788
rect 319713 338738 319779 338741
rect 316572 338736 319779 338738
rect 316572 338728 319718 338736
rect 157198 338678 158871 338680
rect 317094 338680 319718 338728
rect 319774 338680 319779 338736
rect 317094 338678 319779 338680
rect 158805 338675 158871 338678
rect 319713 338675 319779 338678
rect 336733 338602 336799 338605
rect 336733 338600 340124 338602
rect 336733 338544 336738 338600
rect 336794 338544 340124 338600
rect 336733 338542 340124 338544
rect 336733 338539 336799 338542
rect 583520 338452 584960 338692
rect 337745 337922 337811 337925
rect 337745 337920 340124 337922
rect 337745 337864 337750 337920
rect 337806 337864 340124 337920
rect 337745 337862 340124 337864
rect 337745 337859 337811 337862
rect 156588 337242 157258 337292
rect 158989 337242 159055 337245
rect 156588 337240 159055 337242
rect 156588 337232 158994 337240
rect 157198 337184 158994 337232
rect 159050 337184 159055 337240
rect 316572 337242 317154 337292
rect 319805 337242 319871 337245
rect 316572 337240 319871 337242
rect 316572 337232 319810 337240
rect 157198 337182 159055 337184
rect 317094 337184 319810 337232
rect 319866 337184 319871 337240
rect 317094 337182 319871 337184
rect 158989 337179 159055 337182
rect 319805 337179 319871 337182
rect 337653 337242 337719 337245
rect 337653 337240 340124 337242
rect 337653 337184 337658 337240
rect 337714 337184 340124 337240
rect 337653 337182 340124 337184
rect 337653 337179 337719 337182
rect 337837 336562 337903 336565
rect 337837 336560 340124 336562
rect 337837 336504 337842 336560
rect 337898 336504 340124 336560
rect 337837 336502 340124 336504
rect 337837 336499 337903 336502
rect 156588 336018 157258 336068
rect 158897 336018 158963 336021
rect 156588 336016 158963 336018
rect 156588 336008 158902 336016
rect 157198 335960 158902 336008
rect 158958 335960 158963 336016
rect 316572 336018 317154 336068
rect 319897 336018 319963 336021
rect 316572 336016 319963 336018
rect 316572 336008 319902 336016
rect 157198 335958 158963 335960
rect 317094 335960 319902 336008
rect 319958 335960 319963 336016
rect 317094 335958 319963 335960
rect 158897 335955 158963 335958
rect 319897 335955 319963 335958
rect 337653 336018 337719 336021
rect 337653 336016 340124 336018
rect 337653 335960 337658 336016
rect 337714 335960 340124 336016
rect 337653 335958 340124 335960
rect 337653 335955 337719 335958
rect 337561 335338 337627 335341
rect 337561 335336 340124 335338
rect 337561 335280 337566 335336
rect 337622 335280 340124 335336
rect 337561 335278 340124 335280
rect 337561 335275 337627 335278
rect 482369 334930 482435 334933
rect 479964 334928 482435 334930
rect 479964 334872 482374 334928
rect 482430 334872 482435 334928
rect 479964 334870 482435 334872
rect 482369 334867 482435 334870
rect 337745 334658 337811 334661
rect 337745 334656 340124 334658
rect 337745 334600 337750 334656
rect 337806 334600 340124 334656
rect 337745 334598 340124 334600
rect 337745 334595 337811 334598
rect 337653 333978 337719 333981
rect 337653 333976 340124 333978
rect 337653 333920 337658 333976
rect 337714 333920 340124 333976
rect 337653 333918 340124 333920
rect 337653 333915 337719 333918
rect 337745 333434 337811 333437
rect 337745 333432 340124 333434
rect 337745 333376 337750 333432
rect 337806 333376 340124 333432
rect 337745 333374 340124 333376
rect 337745 333371 337811 333374
rect 337745 332754 337811 332757
rect 337745 332752 340124 332754
rect 337745 332696 337750 332752
rect 337806 332696 340124 332752
rect 337745 332694 340124 332696
rect 337745 332691 337811 332694
rect -960 332196 480 332436
rect 17033 332346 17099 332349
rect 19382 332346 20056 332396
rect 17033 332344 20056 332346
rect 17033 332288 17038 332344
rect 17094 332336 20056 332344
rect 177941 332346 178007 332349
rect 179462 332346 180032 332396
rect 177941 332344 180032 332346
rect 17094 332288 19442 332336
rect 17033 332286 19442 332288
rect 177941 332288 177946 332344
rect 178002 332336 180032 332344
rect 178002 332288 179522 332336
rect 177941 332286 179522 332288
rect 17033 332283 17099 332286
rect 177941 332283 178007 332286
rect 337653 332074 337719 332077
rect 337653 332072 340124 332074
rect 337653 332016 337658 332072
rect 337714 332016 340124 332072
rect 337653 332014 340124 332016
rect 337653 332011 337719 332014
rect 336181 331530 336247 331533
rect 336181 331528 340124 331530
rect 336181 331472 336186 331528
rect 336242 331472 340124 331528
rect 336181 331470 340124 331472
rect 336181 331467 336247 331470
rect 176653 330850 176719 330853
rect 337653 330850 337719 330853
rect 176653 330848 179522 330850
rect 176653 330792 176658 330848
rect 176714 330792 179522 330848
rect 176653 330790 179522 330792
rect 176653 330787 176719 330790
rect 179462 330764 179522 330790
rect 337653 330848 340124 330850
rect 337653 330792 337658 330848
rect 337714 330792 340124 330848
rect 337653 330790 340124 330792
rect 337653 330787 337719 330790
rect 17861 330714 17927 330717
rect 19382 330714 20056 330764
rect 17861 330712 20056 330714
rect 17861 330656 17866 330712
rect 17922 330704 20056 330712
rect 179462 330704 180032 330764
rect 17922 330656 19442 330704
rect 17861 330654 19442 330656
rect 17861 330651 17927 330654
rect 17033 330442 17099 330445
rect 19382 330442 20056 330492
rect 17033 330440 20056 330442
rect 17033 330384 17038 330440
rect 17094 330432 20056 330440
rect 177113 330442 177179 330445
rect 177941 330442 178007 330445
rect 179462 330442 180032 330492
rect 177113 330440 180032 330442
rect 17094 330384 19442 330432
rect 17033 330382 19442 330384
rect 177113 330384 177118 330440
rect 177174 330384 177946 330440
rect 178002 330432 180032 330440
rect 178002 330384 179522 330432
rect 177113 330382 179522 330384
rect 17033 330379 17099 330382
rect 177113 330379 177179 330382
rect 177941 330379 178007 330382
rect 482277 330306 482343 330309
rect 479964 330304 482343 330306
rect 479964 330248 482282 330304
rect 482338 330248 482343 330304
rect 479964 330246 482343 330248
rect 482277 330243 482343 330246
rect 337745 330170 337811 330173
rect 337745 330168 340124 330170
rect 337745 330112 337750 330168
rect 337806 330112 340124 330168
rect 337745 330110 340124 330112
rect 337745 330107 337811 330110
rect 337653 329490 337719 329493
rect 337653 329488 340124 329490
rect 337653 329432 337658 329488
rect 337714 329432 340124 329488
rect 337653 329430 340124 329432
rect 337653 329427 337719 329430
rect 337653 328946 337719 328949
rect 337653 328944 340124 328946
rect 337653 328888 337658 328944
rect 337714 328888 340124 328944
rect 337653 328886 340124 328888
rect 337653 328883 337719 328886
rect 337561 328266 337627 328269
rect 337561 328264 340124 328266
rect 337561 328208 337566 328264
rect 337622 328208 340124 328264
rect 337561 328206 340124 328208
rect 337561 328203 337627 328206
rect 337101 327586 337167 327589
rect 337101 327584 340124 327586
rect 337101 327528 337106 327584
rect 337162 327528 340124 327584
rect 337101 327526 340124 327528
rect 337101 327523 337167 327526
rect 337653 327042 337719 327045
rect 337653 327040 340124 327042
rect 337653 326984 337658 327040
rect 337714 326984 340124 327040
rect 337653 326982 340124 326984
rect 337653 326979 337719 326982
rect 337653 326362 337719 326365
rect 337653 326360 340124 326362
rect 337653 326304 337658 326360
rect 337714 326304 340124 326360
rect 337653 326302 340124 326304
rect 337653 326299 337719 326302
rect 337561 325682 337627 325685
rect 482369 325682 482435 325685
rect 337561 325680 340124 325682
rect 337561 325624 337566 325680
rect 337622 325624 340124 325680
rect 337561 325622 340124 325624
rect 479964 325680 482435 325682
rect 479964 325624 482374 325680
rect 482430 325624 482435 325680
rect 479964 325622 482435 325624
rect 337561 325619 337627 325622
rect 482369 325619 482435 325622
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 337653 325002 337719 325005
rect 337653 325000 340124 325002
rect 337653 324944 337658 325000
rect 337714 324944 340124 325000
rect 337653 324942 340124 324944
rect 337653 324939 337719 324942
rect 337745 324458 337811 324461
rect 337745 324456 340124 324458
rect 337745 324400 337750 324456
rect 337806 324400 340124 324456
rect 337745 324398 340124 324400
rect 337745 324395 337811 324398
rect 337653 323778 337719 323781
rect 337653 323776 340124 323778
rect 337653 323720 337658 323776
rect 337714 323720 340124 323776
rect 337653 323718 340124 323720
rect 337653 323715 337719 323718
rect 337469 323098 337535 323101
rect 337469 323096 340124 323098
rect 337469 323040 337474 323096
rect 337530 323040 340124 323096
rect 337469 323038 340124 323040
rect 337469 323035 337535 323038
rect 337745 322554 337811 322557
rect 337745 322552 340124 322554
rect 337745 322496 337750 322552
rect 337806 322496 340124 322552
rect 337745 322494 340124 322496
rect 337745 322491 337811 322494
rect 143349 322012 143415 322013
rect 143349 322008 143358 322012
rect 143422 322010 143428 322012
rect 223481 322010 223547 322013
rect 228633 322012 228699 322013
rect 226926 322010 226932 322012
rect 143349 321952 143354 322008
rect 143349 321948 143358 321952
rect 143422 321950 143506 322010
rect 223481 322008 226932 322010
rect 223481 321952 223486 322008
rect 223542 321952 226932 322008
rect 223481 321950 226932 321952
rect 143422 321948 143428 321950
rect 143349 321947 143415 321948
rect 223481 321947 223547 321950
rect 226926 321948 226932 321950
rect 226996 322010 227002 322012
rect 227600 322010 227606 322012
rect 226996 321950 227606 322010
rect 226996 321948 227002 321950
rect 227600 321948 227606 321950
rect 227670 321948 227676 322012
rect 228633 322008 228694 322012
rect 228633 321952 228638 322008
rect 228633 321948 228694 321952
rect 228758 322010 228764 322012
rect 228758 321950 228790 322010
rect 228758 321948 228764 321950
rect 228633 321947 228699 321948
rect 68686 321812 68692 321876
rect 68756 321874 68762 321876
rect 179638 321874 179644 321876
rect 68756 321814 179644 321874
rect 68756 321812 68762 321814
rect 179638 321812 179644 321814
rect 179708 321874 179714 321876
rect 179781 321874 179847 321877
rect 179708 321872 179847 321874
rect 179708 321816 179786 321872
rect 179842 321816 179847 321872
rect 179708 321814 179847 321816
rect 179708 321812 179714 321814
rect 179781 321811 179847 321814
rect 337653 321874 337719 321877
rect 337653 321872 340124 321874
rect 337653 321816 337658 321872
rect 337714 321816 340124 321872
rect 337653 321814 340124 321816
rect 337653 321811 337719 321814
rect 179413 321740 179479 321741
rect 226333 321740 226399 321741
rect 66478 321676 66484 321740
rect 66548 321738 66554 321740
rect 179413 321738 179460 321740
rect 66548 321736 179460 321738
rect 179524 321738 179530 321740
rect 226333 321738 226380 321740
rect 66548 321680 179418 321736
rect 66548 321678 179460 321680
rect 66548 321676 66554 321678
rect 179413 321676 179460 321678
rect 179524 321678 179606 321738
rect 226288 321736 226380 321738
rect 226288 321680 226338 321736
rect 226288 321678 226380 321680
rect 179524 321676 179530 321678
rect 226333 321676 226380 321678
rect 226444 321676 226450 321740
rect 179413 321675 179479 321676
rect 226333 321675 226399 321676
rect 62757 321604 62823 321605
rect 63861 321604 63927 321605
rect 67633 321604 67699 321605
rect 62757 321600 62804 321604
rect 62868 321602 62874 321604
rect 62757 321544 62762 321600
rect 62757 321540 62804 321544
rect 62868 321542 62914 321602
rect 63861 321600 63908 321604
rect 63972 321602 63978 321604
rect 67582 321602 67588 321604
rect 63861 321544 63866 321600
rect 62868 321540 62874 321542
rect 63861 321540 63908 321544
rect 63972 321542 64018 321602
rect 67506 321542 67588 321602
rect 67652 321602 67699 321604
rect 179505 321602 179571 321605
rect 180006 321602 180012 321604
rect 67652 321600 180012 321602
rect 67694 321544 179510 321600
rect 179566 321544 180012 321600
rect 63972 321540 63978 321542
rect 67582 321540 67588 321542
rect 67652 321542 180012 321544
rect 67652 321540 67699 321542
rect 62757 321539 62823 321540
rect 63861 321539 63927 321540
rect 67633 321539 67699 321540
rect 179505 321539 179571 321542
rect 180006 321540 180012 321542
rect 180076 321540 180082 321604
rect 19006 321404 19012 321468
rect 19076 321466 19082 321468
rect 58198 321466 58204 321468
rect 19076 321406 58204 321466
rect 19076 321404 19082 321406
rect 58198 321404 58204 321406
rect 58268 321466 58274 321468
rect 178953 321466 179019 321469
rect 180149 321466 180215 321469
rect 58268 321464 180215 321466
rect 58268 321408 178958 321464
rect 179014 321408 180154 321464
rect 180210 321408 180215 321464
rect 58268 321406 180215 321408
rect 58268 321404 58274 321406
rect 178953 321403 179019 321406
rect 180149 321403 180215 321406
rect 219198 321404 219204 321468
rect 219268 321466 219274 321468
rect 219433 321466 219499 321469
rect 219268 321464 219499 321466
rect 219268 321408 219438 321464
rect 219494 321408 219499 321464
rect 219268 321406 219499 321408
rect 219268 321404 219274 321406
rect 219433 321403 219499 321406
rect 220445 321466 220511 321469
rect 220670 321466 220676 321468
rect 220445 321464 220676 321466
rect 220445 321408 220450 321464
rect 220506 321408 220676 321464
rect 220445 321406 220676 321408
rect 220445 321403 220511 321406
rect 220670 321404 220676 321406
rect 220740 321404 220746 321468
rect 19190 321268 19196 321332
rect 19260 321330 19266 321332
rect 56910 321330 56916 321332
rect 19260 321270 56916 321330
rect 19260 321268 19266 321270
rect 56910 321268 56916 321270
rect 56980 321330 56986 321332
rect 178125 321330 178191 321333
rect 56980 321328 178191 321330
rect 56980 321272 178130 321328
rect 178186 321272 178191 321328
rect 56980 321270 178191 321272
rect 56980 321268 56986 321270
rect 178125 321267 178191 321270
rect 19425 321194 19491 321197
rect 54518 321194 54524 321196
rect 19425 321192 54524 321194
rect 19425 321136 19430 321192
rect 19486 321136 54524 321192
rect 19425 321134 54524 321136
rect 19425 321131 19491 321134
rect 54518 321132 54524 321134
rect 54588 321194 54594 321196
rect 179505 321194 179571 321197
rect 54588 321192 179571 321194
rect 54588 321136 179510 321192
rect 179566 321136 179571 321192
rect 54588 321134 179571 321136
rect 54588 321132 54594 321134
rect 179505 321131 179571 321134
rect 337653 321194 337719 321197
rect 337653 321192 340124 321194
rect 337653 321136 337658 321192
rect 337714 321136 340124 321192
rect 337653 321134 340124 321136
rect 337653 321131 337719 321134
rect 3417 321058 3483 321061
rect 321185 321058 321251 321061
rect 3417 321056 321251 321058
rect 3417 321000 3422 321056
rect 3478 321000 321190 321056
rect 321246 321000 321251 321056
rect 3417 320998 321251 321000
rect 3417 320995 3483 320998
rect 321185 320995 321251 320998
rect 3785 320922 3851 320925
rect 322473 320922 322539 320925
rect 482277 320922 482343 320925
rect 3785 320920 322539 320922
rect 3785 320864 3790 320920
rect 3846 320864 322478 320920
rect 322534 320864 322539 320920
rect 3785 320862 322539 320864
rect 479964 320920 482343 320922
rect 479964 320864 482282 320920
rect 482338 320864 482343 320920
rect 479964 320862 482343 320864
rect 3785 320859 3851 320862
rect 322473 320859 322539 320862
rect 482277 320859 482343 320862
rect 3601 320786 3667 320789
rect 328085 320786 328151 320789
rect 3601 320784 328151 320786
rect 3601 320728 3606 320784
rect 3662 320728 328090 320784
rect 328146 320728 328151 320784
rect 3601 320726 328151 320728
rect 3601 320723 3667 320726
rect 328085 320723 328151 320726
rect 19374 320588 19380 320652
rect 19444 320650 19450 320652
rect 61694 320650 61700 320652
rect 19444 320590 61700 320650
rect 19444 320588 19450 320590
rect 61694 320588 61700 320590
rect 61764 320650 61770 320652
rect 178033 320650 178099 320653
rect 61764 320648 178099 320650
rect 61764 320592 178038 320648
rect 178094 320592 178099 320648
rect 61764 320590 178099 320592
rect 61764 320588 61770 320590
rect 178033 320587 178099 320590
rect 207289 320650 207355 320653
rect 221825 320652 221891 320653
rect 207606 320650 207612 320652
rect 207289 320648 207612 320650
rect 207289 320592 207294 320648
rect 207350 320592 207612 320648
rect 207289 320590 207612 320592
rect 207289 320587 207355 320590
rect 207606 320588 207612 320590
rect 207676 320588 207682 320652
rect 221774 320650 221780 320652
rect 221734 320590 221780 320650
rect 221844 320648 221891 320652
rect 221886 320592 221891 320648
rect 221774 320588 221780 320590
rect 221844 320588 221891 320592
rect 221825 320587 221891 320588
rect 20662 320452 20668 320516
rect 20732 320514 20738 320516
rect 67633 320514 67699 320517
rect 74625 320516 74691 320517
rect 143257 320516 143323 320517
rect 74574 320514 74580 320516
rect 20732 320512 67699 320514
rect 20732 320456 67638 320512
rect 67694 320456 67699 320512
rect 20732 320454 67699 320456
rect 74534 320454 74580 320514
rect 74644 320512 74691 320516
rect 143206 320514 143212 320516
rect 74686 320456 74691 320512
rect 20732 320452 20738 320454
rect 67633 320451 67699 320454
rect 74574 320452 74580 320454
rect 74644 320452 74691 320456
rect 143166 320454 143212 320514
rect 143276 320512 143323 320516
rect 143318 320456 143323 320512
rect 143206 320452 143212 320454
rect 143276 320452 143323 320456
rect 74625 320451 74691 320452
rect 143257 320451 143323 320452
rect 336917 320514 336983 320517
rect 336917 320512 340124 320514
rect 336917 320456 336922 320512
rect 336978 320456 340124 320512
rect 336917 320454 340124 320456
rect 336917 320451 336983 320454
rect 178585 320244 178651 320245
rect 178769 320244 178835 320245
rect 43110 320242 43116 320244
rect 42750 320182 43116 320242
rect 42750 320106 42810 320182
rect 43110 320180 43116 320182
rect 43180 320242 43186 320244
rect 178534 320242 178540 320244
rect 43180 320182 178540 320242
rect 178604 320240 178651 320244
rect 178646 320184 178651 320240
rect 43180 320180 43186 320182
rect 178534 320180 178540 320182
rect 178604 320180 178651 320184
rect 178718 320180 178724 320244
rect 178788 320242 178835 320244
rect 179505 320242 179571 320245
rect 179822 320242 179828 320244
rect 178788 320240 178880 320242
rect 178830 320184 178880 320240
rect 178788 320182 178880 320184
rect 179505 320240 179828 320242
rect 179505 320184 179510 320240
rect 179566 320184 179828 320240
rect 179505 320182 179828 320184
rect 178788 320180 178835 320182
rect 178585 320179 178651 320180
rect 178769 320179 178835 320180
rect 179505 320179 179571 320182
rect 179822 320180 179828 320182
rect 179892 320180 179898 320244
rect 26190 320046 42810 320106
rect 44173 320108 44239 320109
rect 45001 320108 45067 320109
rect 50153 320108 50219 320109
rect 51257 320108 51323 320109
rect 52361 320108 52427 320109
rect 53465 320108 53531 320109
rect 59353 320108 59419 320109
rect 44173 320104 44220 320108
rect 44284 320106 44290 320108
rect 44950 320106 44956 320108
rect 44173 320048 44178 320104
rect 18822 319772 18828 319836
rect 18892 319834 18898 319836
rect 26190 319834 26250 320046
rect 44173 320044 44220 320048
rect 44284 320046 44330 320106
rect 44910 320046 44956 320106
rect 45020 320104 45067 320108
rect 50102 320106 50108 320108
rect 45062 320048 45067 320104
rect 44284 320044 44290 320046
rect 44950 320044 44956 320046
rect 45020 320044 45067 320048
rect 50062 320046 50108 320106
rect 50172 320104 50219 320108
rect 51206 320106 51212 320108
rect 50214 320048 50219 320104
rect 50102 320044 50108 320046
rect 50172 320044 50219 320048
rect 51166 320046 51212 320106
rect 51276 320104 51323 320108
rect 52310 320106 52316 320108
rect 51318 320048 51323 320104
rect 51206 320044 51212 320046
rect 51276 320044 51323 320048
rect 52270 320046 52316 320106
rect 52380 320104 52427 320108
rect 53414 320106 53420 320108
rect 52422 320048 52427 320104
rect 52310 320044 52316 320046
rect 52380 320044 52427 320048
rect 53374 320046 53420 320106
rect 53484 320104 53531 320108
rect 59302 320106 59308 320108
rect 53526 320048 53531 320104
rect 53414 320044 53420 320046
rect 53484 320044 53531 320048
rect 59226 320046 59308 320106
rect 59372 320106 59419 320108
rect 60641 320106 60707 320109
rect 59372 320104 60707 320106
rect 59414 320048 60646 320104
rect 60702 320048 60707 320104
rect 59302 320044 59308 320046
rect 59372 320046 60707 320048
rect 59372 320044 59419 320046
rect 44173 320043 44239 320044
rect 45001 320043 45067 320044
rect 50153 320043 50219 320044
rect 51257 320043 51323 320044
rect 52361 320043 52427 320044
rect 53465 320043 53531 320044
rect 59353 320043 59419 320044
rect 60641 320043 60707 320046
rect 65333 320108 65399 320109
rect 68645 320108 68711 320109
rect 71129 320108 71195 320109
rect 65333 320104 65380 320108
rect 65444 320106 65450 320108
rect 65333 320048 65338 320104
rect 65333 320044 65380 320048
rect 65444 320046 65490 320106
rect 68645 320104 68692 320108
rect 68756 320106 68762 320108
rect 71078 320106 71084 320108
rect 68645 320048 68650 320104
rect 65444 320044 65450 320046
rect 68645 320044 68692 320048
rect 68756 320046 68802 320106
rect 71038 320046 71084 320106
rect 71148 320104 71195 320108
rect 71190 320048 71195 320104
rect 68756 320044 68762 320046
rect 71078 320044 71084 320046
rect 71148 320044 71195 320048
rect 65333 320043 65399 320044
rect 68645 320043 68711 320044
rect 71129 320043 71195 320044
rect 72141 320108 72207 320109
rect 73337 320108 73403 320109
rect 75729 320108 75795 320109
rect 79225 320108 79291 320109
rect 72141 320104 72188 320108
rect 72252 320106 72258 320108
rect 73286 320106 73292 320108
rect 72141 320048 72146 320104
rect 72141 320044 72188 320048
rect 72252 320046 72298 320106
rect 73246 320046 73292 320106
rect 73356 320104 73403 320108
rect 75678 320106 75684 320108
rect 73398 320048 73403 320104
rect 72252 320044 72258 320046
rect 73286 320044 73292 320046
rect 73356 320044 73403 320048
rect 75638 320046 75684 320106
rect 75748 320104 75795 320108
rect 79174 320106 79180 320108
rect 75790 320048 75795 320104
rect 75678 320044 75684 320046
rect 75748 320044 75795 320048
rect 79134 320046 79180 320106
rect 79244 320104 79291 320108
rect 79286 320048 79291 320104
rect 79174 320044 79180 320046
rect 79244 320044 79291 320048
rect 200614 320044 200620 320108
rect 200684 320106 200690 320108
rect 200757 320106 200823 320109
rect 203149 320108 203215 320109
rect 203149 320106 203196 320108
rect 200684 320104 200823 320106
rect 200684 320048 200762 320104
rect 200818 320048 200823 320104
rect 200684 320046 200823 320048
rect 203068 320104 203196 320106
rect 203260 320106 203266 320108
rect 203793 320106 203859 320109
rect 204345 320108 204411 320109
rect 204294 320106 204300 320108
rect 203260 320104 203859 320106
rect 203068 320048 203154 320104
rect 203260 320048 203798 320104
rect 203854 320048 203859 320104
rect 203068 320046 203196 320048
rect 200684 320044 200690 320046
rect 72141 320043 72207 320044
rect 73337 320043 73403 320044
rect 75729 320043 75795 320044
rect 79225 320043 79291 320044
rect 200757 320043 200823 320046
rect 203149 320044 203196 320046
rect 203260 320046 203859 320048
rect 204254 320046 204300 320106
rect 204364 320104 204411 320108
rect 204406 320048 204411 320104
rect 203260 320044 203266 320046
rect 203149 320043 203215 320044
rect 203793 320043 203859 320046
rect 204294 320044 204300 320046
rect 204364 320044 204411 320048
rect 211654 320044 211660 320108
rect 211724 320106 211730 320108
rect 211797 320106 211863 320109
rect 211724 320104 211863 320106
rect 211724 320048 211802 320104
rect 211858 320048 211863 320104
rect 211724 320046 211863 320048
rect 211724 320044 211730 320046
rect 204345 320043 204411 320044
rect 211797 320043 211863 320046
rect 223982 320044 223988 320108
rect 224052 320106 224058 320108
rect 224125 320106 224191 320109
rect 224052 320104 224191 320106
rect 224052 320048 224130 320104
rect 224186 320048 224191 320104
rect 224052 320046 224191 320048
rect 224052 320044 224058 320046
rect 224125 320043 224191 320046
rect 226374 320044 226380 320108
rect 226444 320106 226450 320108
rect 227529 320106 227595 320109
rect 231209 320108 231275 320109
rect 231158 320106 231164 320108
rect 226444 320104 227595 320106
rect 226444 320048 227534 320104
rect 227590 320048 227595 320104
rect 226444 320046 227595 320048
rect 231118 320046 231164 320106
rect 231228 320104 231275 320108
rect 231270 320048 231275 320104
rect 226444 320044 226450 320046
rect 227529 320043 227595 320046
rect 231158 320044 231164 320046
rect 231228 320044 231275 320048
rect 231209 320043 231275 320044
rect 36077 319972 36143 319973
rect 39573 319972 39639 319973
rect 36077 319968 36124 319972
rect 36188 319970 36194 319972
rect 36077 319912 36082 319968
rect 36077 319908 36124 319912
rect 36188 319910 36234 319970
rect 39573 319968 39620 319972
rect 39684 319970 39690 319972
rect 59905 319970 59971 319973
rect 60590 319970 60596 319972
rect 39573 319912 39578 319968
rect 36188 319908 36194 319910
rect 39573 319908 39620 319912
rect 39684 319910 39730 319970
rect 59905 319968 60596 319970
rect 59905 319912 59910 319968
rect 59966 319912 60596 319968
rect 59905 319910 60596 319912
rect 39684 319908 39690 319910
rect 36077 319907 36143 319908
rect 39573 319907 39639 319908
rect 59905 319907 59971 319910
rect 60590 319908 60596 319910
rect 60660 319970 60666 319972
rect 60825 319970 60891 319973
rect 66437 319972 66503 319973
rect 66437 319970 66484 319972
rect 60660 319968 60891 319970
rect 60660 319912 60830 319968
rect 60886 319912 60891 319968
rect 60660 319910 60891 319912
rect 66392 319968 66484 319970
rect 66392 319912 66442 319968
rect 66392 319910 66484 319912
rect 60660 319908 60666 319910
rect 60825 319907 60891 319910
rect 66437 319908 66484 319910
rect 66548 319908 66554 319972
rect 214598 319908 214604 319972
rect 214668 319970 214674 319972
rect 215109 319970 215175 319973
rect 226977 319972 227043 319973
rect 214668 319968 215175 319970
rect 214668 319912 215114 319968
rect 215170 319912 215175 319968
rect 214668 319910 215175 319912
rect 214668 319908 214674 319910
rect 66437 319907 66503 319908
rect 215109 319907 215175 319910
rect 226926 319908 226932 319972
rect 226996 319970 227043 319972
rect 229553 319970 229619 319973
rect 229686 319970 229692 319972
rect 226996 319968 227088 319970
rect 227038 319912 227088 319968
rect 226996 319910 227088 319912
rect 229553 319968 229692 319970
rect 229553 319912 229558 319968
rect 229614 319912 229692 319968
rect 229553 319910 229692 319912
rect 226996 319908 227043 319910
rect 226977 319907 227043 319908
rect 229553 319907 229619 319910
rect 229686 319908 229692 319910
rect 229756 319908 229762 319972
rect 337745 319970 337811 319973
rect 337745 319968 340124 319970
rect 337745 319912 337750 319968
rect 337806 319912 340124 319968
rect 337745 319910 340124 319912
rect 337745 319907 337811 319910
rect 18892 319774 26250 319834
rect 18892 319772 18898 319774
rect 209998 319772 210004 319836
rect 210068 319834 210074 319836
rect 210417 319834 210483 319837
rect 210068 319832 210483 319834
rect 210068 319776 210422 319832
rect 210478 319776 210483 319832
rect 210068 319774 210483 319776
rect 210068 319772 210074 319774
rect 210417 319771 210483 319774
rect 18689 319698 18755 319701
rect 55622 319698 55628 319700
rect 18689 319696 55628 319698
rect 18689 319640 18694 319696
rect 18750 319640 55628 319696
rect 18689 319638 55628 319640
rect 18689 319635 18755 319638
rect 55622 319636 55628 319638
rect 55692 319698 55698 319700
rect 56501 319698 56567 319701
rect 55692 319696 56567 319698
rect 55692 319640 56506 319696
rect 56562 319640 56567 319696
rect 55692 319638 56567 319640
rect 55692 319636 55698 319638
rect 56501 319635 56567 319638
rect 78254 319636 78260 319700
rect 78324 319698 78330 319700
rect 78673 319698 78739 319701
rect 78324 319696 78739 319698
rect 78324 319640 78678 319696
rect 78734 319640 78739 319696
rect 78324 319638 78739 319640
rect 78324 319636 78330 319638
rect 78673 319635 78739 319638
rect 215886 319636 215892 319700
rect 215956 319698 215962 319700
rect 216397 319698 216463 319701
rect 215956 319696 216463 319698
rect 215956 319640 216402 319696
rect 216458 319640 216463 319696
rect 215956 319638 216463 319640
rect 215956 319636 215962 319638
rect 216397 319635 216463 319638
rect 216673 319698 216739 319701
rect 216990 319698 216996 319700
rect 216673 319696 216996 319698
rect 216673 319640 216678 319696
rect 216734 319640 216996 319696
rect 216673 319638 216996 319640
rect 216673 319635 216739 319638
rect 216990 319636 216996 319638
rect 217060 319698 217066 319700
rect 217869 319698 217935 319701
rect 217060 319696 217935 319698
rect 217060 319640 217874 319696
rect 217930 319640 217935 319696
rect 217060 319638 217935 319640
rect 217060 319636 217066 319638
rect 217869 319635 217935 319638
rect 218053 319698 218119 319701
rect 218646 319698 218652 319700
rect 218053 319696 218652 319698
rect 218053 319640 218058 319696
rect 218114 319640 218652 319696
rect 218053 319638 218652 319640
rect 218053 319635 218119 319638
rect 218646 319636 218652 319638
rect 218716 319698 218722 319700
rect 219249 319698 219315 319701
rect 218716 319696 219315 319698
rect 218716 319640 219254 319696
rect 219310 319640 219315 319696
rect 218716 319638 219315 319640
rect 218716 319636 218722 319638
rect 219249 319635 219315 319638
rect 231853 319698 231919 319701
rect 232262 319698 232268 319700
rect 231853 319696 232268 319698
rect 231853 319640 231858 319696
rect 231914 319640 232268 319696
rect 231853 319638 232268 319640
rect 231853 319635 231919 319638
rect 232262 319636 232268 319638
rect 232332 319698 232338 319700
rect 232497 319698 232563 319701
rect 232332 319696 232563 319698
rect 232332 319640 232502 319696
rect 232558 319640 232563 319696
rect 232332 319638 232563 319640
rect 232332 319636 232338 319638
rect 232497 319635 232563 319638
rect 18638 319500 18644 319564
rect 18708 319562 18714 319564
rect 48630 319562 48636 319564
rect 18708 319502 48636 319562
rect 18708 319500 18714 319502
rect 48630 319500 48636 319502
rect 48700 319562 48706 319564
rect 179270 319562 179276 319564
rect 48700 319502 179276 319562
rect 48700 319500 48706 319502
rect 179270 319500 179276 319502
rect 179340 319562 179346 319564
rect 236637 319562 236703 319565
rect 236862 319562 236868 319564
rect 179340 319502 180810 319562
rect 179340 319500 179346 319502
rect -960 319140 480 319380
rect 19558 319364 19564 319428
rect 19628 319426 19634 319428
rect 47526 319426 47532 319428
rect 19628 319366 47532 319426
rect 19628 319364 19634 319366
rect 47526 319364 47532 319366
rect 47596 319426 47602 319428
rect 178033 319426 178099 319429
rect 179086 319426 179092 319428
rect 47596 319424 179092 319426
rect 47596 319368 178038 319424
rect 178094 319368 179092 319424
rect 47596 319366 179092 319368
rect 47596 319364 47602 319366
rect 178033 319363 178099 319366
rect 179086 319364 179092 319366
rect 179156 319364 179162 319428
rect 40534 319228 40540 319292
rect 40604 319290 40610 319292
rect 40677 319290 40743 319293
rect 40604 319288 40743 319290
rect 40604 319232 40682 319288
rect 40738 319232 40743 319288
rect 40604 319230 40743 319232
rect 40604 319228 40610 319230
rect 40677 319227 40743 319230
rect 42057 319290 42123 319293
rect 42374 319290 42380 319292
rect 42057 319288 42380 319290
rect 42057 319232 42062 319288
rect 42118 319232 42380 319288
rect 42057 319230 42380 319232
rect 42057 319227 42123 319230
rect 42374 319228 42380 319230
rect 42444 319228 42450 319292
rect 69790 319228 69796 319292
rect 69860 319290 69866 319292
rect 70393 319290 70459 319293
rect 69860 319288 70459 319290
rect 69860 319232 70398 319288
rect 70454 319232 70459 319288
rect 69860 319230 70459 319232
rect 69860 319228 69866 319230
rect 70393 319227 70459 319230
rect 76966 319228 76972 319292
rect 77036 319290 77042 319292
rect 77293 319290 77359 319293
rect 77036 319288 77359 319290
rect 77036 319232 77298 319288
rect 77354 319232 77359 319288
rect 77036 319230 77359 319232
rect 180750 319290 180810 319502
rect 236637 319560 236868 319562
rect 236637 319504 236642 319560
rect 236698 319504 236868 319560
rect 236637 319502 236868 319504
rect 236637 319499 236703 319502
rect 236862 319500 236868 319502
rect 236932 319500 236938 319564
rect 196065 319428 196131 319429
rect 196014 319364 196020 319428
rect 196084 319426 196131 319428
rect 197353 319426 197419 319429
rect 198222 319426 198228 319428
rect 196084 319424 196176 319426
rect 196126 319368 196176 319424
rect 196084 319366 196176 319368
rect 197353 319424 198228 319426
rect 197353 319368 197358 319424
rect 197414 319368 198228 319424
rect 197353 319366 198228 319368
rect 196084 319364 196131 319366
rect 196065 319363 196131 319364
rect 197353 319363 197419 319366
rect 198222 319364 198228 319366
rect 198292 319364 198298 319428
rect 198733 319426 198799 319429
rect 199510 319426 199516 319428
rect 198733 319424 199516 319426
rect 198733 319368 198738 319424
rect 198794 319368 199516 319424
rect 198733 319366 199516 319368
rect 198733 319363 198799 319366
rect 199510 319364 199516 319366
rect 199580 319364 199586 319428
rect 213177 319426 213243 319429
rect 222837 319428 222903 319429
rect 303061 319428 303127 319429
rect 213494 319426 213500 319428
rect 200070 319366 208778 319426
rect 200070 319290 200130 319366
rect 180750 319230 200130 319290
rect 201493 319290 201559 319293
rect 201718 319290 201724 319292
rect 201493 319288 201724 319290
rect 201493 319232 201498 319288
rect 201554 319232 201724 319288
rect 201493 319230 201724 319232
rect 77036 319228 77042 319230
rect 77293 319227 77359 319230
rect 201493 319227 201559 319230
rect 201718 319228 201724 319230
rect 201788 319228 201794 319292
rect 206277 319290 206343 319293
rect 208718 319292 208778 319366
rect 213177 319424 213500 319426
rect 213177 319368 213182 319424
rect 213238 319368 213500 319424
rect 213177 319366 213500 319368
rect 213177 319363 213243 319366
rect 213494 319364 213500 319366
rect 213564 319364 213570 319428
rect 222837 319426 222884 319428
rect 222792 319424 222884 319426
rect 222792 319368 222842 319424
rect 222792 319366 222884 319368
rect 222837 319364 222884 319366
rect 222948 319364 222954 319428
rect 303061 319426 303108 319428
rect 303016 319424 303108 319426
rect 303016 319368 303066 319424
rect 303016 319366 303108 319368
rect 303061 319364 303108 319366
rect 303172 319364 303178 319428
rect 222837 319363 222903 319364
rect 303061 319363 303127 319364
rect 206502 319290 206508 319292
rect 204118 319288 206508 319290
rect 204118 319232 206282 319288
rect 206338 319232 206508 319288
rect 204118 319230 206508 319232
rect 36537 319154 36603 319157
rect 37038 319154 37044 319156
rect 36537 319152 37044 319154
rect 36537 319096 36542 319152
rect 36598 319096 37044 319152
rect 36537 319094 37044 319096
rect 36537 319091 36603 319094
rect 37038 319092 37044 319094
rect 37108 319092 37114 319156
rect 37917 319154 37983 319157
rect 38510 319154 38516 319156
rect 37917 319152 38516 319154
rect 37917 319096 37922 319152
rect 37978 319096 38516 319152
rect 37917 319094 38516 319096
rect 37917 319091 37983 319094
rect 38510 319092 38516 319094
rect 38580 319092 38586 319156
rect 46197 319154 46263 319157
rect 46422 319154 46428 319156
rect 46197 319152 46428 319154
rect 46197 319096 46202 319152
rect 46258 319096 46428 319152
rect 46197 319094 46428 319096
rect 46197 319091 46263 319094
rect 46422 319092 46428 319094
rect 46492 319092 46498 319156
rect 177982 319092 177988 319156
rect 178052 319154 178058 319156
rect 178902 319154 178908 319156
rect 178052 319094 178908 319154
rect 178052 319092 178058 319094
rect 178902 319092 178908 319094
rect 178972 319154 178978 319156
rect 204118 319154 204178 319230
rect 206277 319227 206343 319230
rect 206502 319228 206508 319230
rect 206572 319228 206578 319292
rect 208710 319228 208716 319292
rect 208780 319290 208786 319292
rect 209037 319290 209103 319293
rect 208780 319288 209103 319290
rect 208780 319232 209042 319288
rect 209098 319232 209103 319288
rect 208780 319230 209103 319232
rect 208780 319228 208786 319230
rect 209037 319227 209103 319230
rect 224902 319228 224908 319292
rect 224972 319290 224978 319292
rect 225597 319290 225663 319293
rect 224972 319288 225663 319290
rect 224972 319232 225602 319288
rect 225658 319232 225663 319288
rect 224972 319230 225663 319232
rect 224972 319228 224978 319230
rect 225597 319227 225663 319230
rect 234061 319290 234127 319293
rect 234286 319290 234292 319292
rect 234061 319288 234292 319290
rect 234061 319232 234066 319288
rect 234122 319232 234292 319288
rect 234061 319230 234292 319232
rect 234061 319227 234127 319230
rect 234286 319228 234292 319230
rect 234356 319228 234362 319292
rect 235257 319290 235323 319293
rect 235574 319290 235580 319292
rect 235257 319288 235580 319290
rect 235257 319232 235262 319288
rect 235318 319232 235580 319288
rect 235257 319230 235580 319232
rect 235257 319227 235323 319230
rect 235574 319228 235580 319230
rect 235644 319228 235650 319292
rect 302877 319290 302943 319293
rect 303470 319290 303476 319292
rect 302877 319288 303476 319290
rect 302877 319232 302882 319288
rect 302938 319232 303476 319288
rect 302877 319230 303476 319232
rect 302877 319227 302943 319230
rect 303470 319228 303476 319230
rect 303540 319228 303546 319292
rect 337653 319290 337719 319293
rect 337653 319288 340124 319290
rect 337653 319232 337658 319288
rect 337714 319232 340124 319288
rect 337653 319230 340124 319232
rect 337653 319227 337719 319230
rect 178972 319094 204178 319154
rect 204253 319154 204319 319157
rect 205398 319154 205404 319156
rect 204253 319152 205404 319154
rect 204253 319096 204258 319152
rect 204314 319096 205404 319152
rect 204253 319094 205404 319096
rect 178972 319092 178978 319094
rect 204253 319091 204319 319094
rect 205398 319092 205404 319094
rect 205468 319092 205474 319156
rect 211337 319154 211403 319157
rect 211981 319154 212047 319157
rect 238017 319156 238083 319157
rect 212390 319154 212396 319156
rect 211337 319152 212396 319154
rect 211337 319096 211342 319152
rect 211398 319096 211986 319152
rect 212042 319096 212396 319152
rect 211337 319094 212396 319096
rect 211337 319091 211403 319094
rect 211981 319091 212047 319094
rect 212390 319092 212396 319094
rect 212460 319092 212466 319156
rect 237966 319092 237972 319156
rect 238036 319154 238083 319156
rect 238036 319152 238128 319154
rect 238078 319096 238128 319152
rect 238036 319094 238128 319096
rect 238036 319092 238083 319094
rect 238017 319091 238083 319092
rect 157333 319018 157399 319021
rect 239070 319018 239076 319020
rect 157333 319016 239076 319018
rect 157333 318960 157338 319016
rect 157394 318960 239076 319016
rect 157333 318958 239076 318960
rect 157333 318955 157399 318958
rect 239070 318956 239076 318958
rect 239140 319018 239146 319020
rect 239397 319018 239463 319021
rect 239140 319016 239463 319018
rect 239140 318960 239402 319016
rect 239458 318960 239463 319016
rect 239140 318958 239463 318960
rect 239140 318956 239146 318958
rect 239397 318955 239463 318958
rect 46197 318882 46263 318885
rect 180517 318884 180583 318885
rect 177982 318882 177988 318884
rect 46197 318880 177988 318882
rect 46197 318824 46202 318880
rect 46258 318824 177988 318880
rect 46197 318822 177988 318824
rect 46197 318819 46263 318822
rect 177982 318820 177988 318822
rect 178052 318820 178058 318884
rect 180517 318880 180564 318884
rect 180628 318882 180634 318884
rect 195973 318882 196039 318885
rect 197118 318882 197124 318884
rect 180517 318824 180522 318880
rect 180517 318820 180564 318824
rect 180628 318822 180674 318882
rect 195973 318880 197124 318882
rect 195973 318824 195978 318880
rect 196034 318824 197124 318880
rect 195973 318822 197124 318824
rect 180628 318820 180634 318822
rect 180517 318819 180583 318820
rect 195973 318819 196039 318822
rect 197118 318820 197124 318822
rect 197188 318820 197194 318884
rect 233366 318820 233372 318884
rect 233436 318882 233442 318884
rect 233877 318882 233943 318885
rect 233436 318880 233943 318882
rect 233436 318824 233882 318880
rect 233938 318824 233943 318880
rect 233436 318822 233943 318824
rect 233436 318820 233442 318822
rect 233877 318819 233943 318822
rect 336917 318610 336983 318613
rect 336917 318608 340124 318610
rect 336917 318552 336922 318608
rect 336978 318552 340124 318608
rect 336917 318550 340124 318552
rect 336917 318547 336983 318550
rect 337653 317930 337719 317933
rect 337653 317928 340124 317930
rect 337653 317872 337658 317928
rect 337714 317872 340124 317928
rect 337653 317870 340124 317872
rect 337653 317867 337719 317870
rect 337561 317386 337627 317389
rect 337561 317384 340124 317386
rect 337561 317328 337566 317384
rect 337622 317328 340124 317384
rect 337561 317326 340124 317328
rect 337561 317323 337627 317326
rect 337653 316706 337719 316709
rect 337653 316704 340124 316706
rect 337653 316648 337658 316704
rect 337714 316648 340124 316704
rect 337653 316646 340124 316648
rect 337653 316643 337719 316646
rect 19558 316236 19564 316300
rect 19628 316298 19634 316300
rect 19793 316298 19859 316301
rect 482001 316298 482067 316301
rect 19628 316296 19859 316298
rect 19628 316240 19798 316296
rect 19854 316240 19859 316296
rect 19628 316238 19859 316240
rect 479964 316296 482067 316298
rect 479964 316240 482006 316296
rect 482062 316240 482067 316296
rect 479964 316238 482067 316240
rect 19628 316236 19634 316238
rect 19793 316235 19859 316238
rect 482001 316235 482067 316238
rect 19425 316162 19491 316165
rect 19558 316162 19564 316164
rect 19425 316160 19564 316162
rect 19425 316104 19430 316160
rect 19486 316104 19564 316160
rect 19425 316102 19564 316104
rect 19425 316099 19491 316102
rect 19558 316100 19564 316102
rect 19628 316100 19634 316164
rect 19374 315964 19380 316028
rect 19444 316026 19450 316028
rect 337745 316026 337811 316029
rect 19444 315966 20730 316026
rect 19444 315964 19450 315966
rect 19374 315828 19380 315892
rect 19444 315890 19450 315892
rect 19793 315890 19859 315893
rect 20670 315892 20730 315966
rect 337745 316024 340124 316026
rect 337745 315968 337750 316024
rect 337806 315968 340124 316024
rect 337745 315966 340124 315968
rect 337745 315963 337811 315966
rect 19444 315888 19859 315890
rect 19444 315832 19798 315888
rect 19854 315832 19859 315888
rect 19444 315830 19859 315832
rect 19444 315828 19450 315830
rect 19793 315827 19859 315830
rect 20662 315828 20668 315892
rect 20732 315828 20738 315892
rect 337653 315482 337719 315485
rect 337653 315480 340124 315482
rect 337653 315424 337658 315480
rect 337714 315424 340124 315480
rect 337653 315422 340124 315424
rect 337653 315419 337719 315422
rect 337653 314802 337719 314805
rect 337653 314800 340124 314802
rect 337653 314744 337658 314800
rect 337714 314744 340124 314800
rect 337653 314742 340124 314744
rect 337653 314739 337719 314742
rect 337653 314122 337719 314125
rect 337653 314120 340124 314122
rect 337653 314064 337658 314120
rect 337714 314064 340124 314120
rect 337653 314062 340124 314064
rect 337653 314059 337719 314062
rect 337653 313442 337719 313445
rect 337653 313440 340124 313442
rect 337653 313384 337658 313440
rect 337714 313384 340124 313440
rect 337653 313382 340124 313384
rect 337653 313379 337719 313382
rect 337745 312898 337811 312901
rect 337745 312896 340124 312898
rect 337745 312840 337750 312896
rect 337806 312840 340124 312896
rect 337745 312838 340124 312840
rect 337745 312835 337811 312838
rect 337745 312218 337811 312221
rect 337745 312216 340124 312218
rect 337745 312160 337750 312216
rect 337806 312160 340124 312216
rect 337745 312158 340124 312160
rect 337745 312155 337811 312158
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 574940 312022 584960 312082
rect 574940 312020 574946 312022
rect 583520 311932 584960 312022
rect 482093 311674 482159 311677
rect 479964 311672 482159 311674
rect 479964 311616 482098 311672
rect 482154 311616 482159 311672
rect 479964 311614 482159 311616
rect 482093 311611 482159 311614
rect 337653 311538 337719 311541
rect 337653 311536 340124 311538
rect 337653 311480 337658 311536
rect 337714 311480 340124 311536
rect 337653 311478 340124 311480
rect 337653 311475 337719 311478
rect 337653 310994 337719 310997
rect 337653 310992 340124 310994
rect 337653 310936 337658 310992
rect 337714 310936 340124 310992
rect 337653 310934 340124 310936
rect 337653 310931 337719 310934
rect 337101 310314 337167 310317
rect 337101 310312 340124 310314
rect 337101 310256 337106 310312
rect 337162 310256 340124 310312
rect 337101 310254 340124 310256
rect 337101 310251 337167 310254
rect 337653 309634 337719 309637
rect 337653 309632 340124 309634
rect 337653 309576 337658 309632
rect 337714 309576 340124 309632
rect 337653 309574 340124 309576
rect 337653 309571 337719 309574
rect 337101 308954 337167 308957
rect 337101 308952 340124 308954
rect 337101 308896 337106 308952
rect 337162 308896 340124 308952
rect 337101 308894 340124 308896
rect 337101 308891 337167 308894
rect 337653 308410 337719 308413
rect 337653 308408 340124 308410
rect 337653 308352 337658 308408
rect 337714 308352 340124 308408
rect 337653 308350 340124 308352
rect 337653 308347 337719 308350
rect 337377 307730 337443 307733
rect 337377 307728 340124 307730
rect 337377 307672 337382 307728
rect 337438 307672 340124 307728
rect 337377 307670 340124 307672
rect 337377 307667 337443 307670
rect 337653 307050 337719 307053
rect 482185 307050 482251 307053
rect 337653 307048 340124 307050
rect 337653 306992 337658 307048
rect 337714 306992 340124 307048
rect 337653 306990 340124 306992
rect 479964 307048 482251 307050
rect 479964 306992 482190 307048
rect 482246 306992 482251 307048
rect 479964 306990 482251 306992
rect 337653 306987 337719 306990
rect 482185 306987 482251 306990
rect 19374 306580 19380 306644
rect 19444 306642 19450 306644
rect 19793 306642 19859 306645
rect 19444 306640 19859 306642
rect 19444 306584 19798 306640
rect 19854 306584 19859 306640
rect 19444 306582 19859 306584
rect 19444 306580 19450 306582
rect 19793 306579 19859 306582
rect 19374 306444 19380 306508
rect 19444 306506 19450 306508
rect 20846 306506 20852 306508
rect 19444 306446 20852 306506
rect 19444 306444 19450 306446
rect 20846 306444 20852 306446
rect 20916 306444 20922 306508
rect 337745 306506 337811 306509
rect 337745 306504 340124 306506
rect 337745 306448 337750 306504
rect 337806 306448 340124 306504
rect 337745 306446 340124 306448
rect 337745 306443 337811 306446
rect -960 306234 480 306324
rect 19374 306308 19380 306372
rect 19444 306370 19450 306372
rect 20846 306370 20852 306372
rect 19444 306310 20852 306370
rect 19444 306308 19450 306310
rect 20846 306308 20852 306310
rect 20916 306308 20922 306372
rect 3785 306234 3851 306237
rect -960 306232 3851 306234
rect -960 306176 3790 306232
rect 3846 306176 3851 306232
rect -960 306174 3851 306176
rect -960 306084 480 306174
rect 3785 306171 3851 306174
rect 19374 306172 19380 306236
rect 19444 306234 19450 306236
rect 19793 306234 19859 306237
rect 19444 306232 19859 306234
rect 19444 306176 19798 306232
rect 19854 306176 19859 306232
rect 19444 306174 19859 306176
rect 19444 306172 19450 306174
rect 19793 306171 19859 306174
rect 337653 305826 337719 305829
rect 337653 305824 340124 305826
rect 337653 305768 337658 305824
rect 337714 305768 340124 305824
rect 337653 305766 340124 305768
rect 337653 305763 337719 305766
rect 337745 305146 337811 305149
rect 337745 305144 340124 305146
rect 337745 305088 337750 305144
rect 337806 305088 340124 305144
rect 337745 305086 340124 305088
rect 337745 305083 337811 305086
rect 337653 304466 337719 304469
rect 337653 304464 340124 304466
rect 337653 304408 337658 304464
rect 337714 304408 340124 304464
rect 337653 304406 340124 304408
rect 337653 304403 337719 304406
rect 337745 303922 337811 303925
rect 337745 303920 340124 303922
rect 337745 303864 337750 303920
rect 337806 303864 340124 303920
rect 337745 303862 340124 303864
rect 337745 303859 337811 303862
rect 337653 303242 337719 303245
rect 337653 303240 340124 303242
rect 337653 303184 337658 303240
rect 337714 303184 340124 303240
rect 337653 303182 340124 303184
rect 337653 303179 337719 303182
rect 336917 302562 336983 302565
rect 336917 302560 340124 302562
rect 336917 302504 336922 302560
rect 336978 302504 340124 302560
rect 336917 302502 340124 302504
rect 336917 302499 336983 302502
rect 482921 302290 482987 302293
rect 479964 302288 482987 302290
rect 479964 302232 482926 302288
rect 482982 302232 482987 302288
rect 479964 302230 482987 302232
rect 482921 302227 482987 302230
rect 337653 301882 337719 301885
rect 337653 301880 340124 301882
rect 337653 301824 337658 301880
rect 337714 301824 340124 301880
rect 337653 301822 340124 301824
rect 337653 301819 337719 301822
rect 337469 301338 337535 301341
rect 337469 301336 340124 301338
rect 337469 301280 337474 301336
rect 337530 301280 340124 301336
rect 337469 301278 340124 301280
rect 337469 301275 337535 301278
rect 337653 300658 337719 300661
rect 337653 300656 340124 300658
rect 337653 300600 337658 300656
rect 337714 300600 340124 300656
rect 337653 300598 340124 300600
rect 337653 300595 337719 300598
rect 337377 299978 337443 299981
rect 337377 299976 340124 299978
rect 337377 299920 337382 299976
rect 337438 299920 340124 299976
rect 337377 299918 340124 299920
rect 337377 299915 337443 299918
rect 337101 299434 337167 299437
rect 337101 299432 340124 299434
rect 337101 299376 337106 299432
rect 337162 299376 340124 299432
rect 337101 299374 340124 299376
rect 337101 299371 337167 299374
rect 337285 298754 337351 298757
rect 337285 298752 340124 298754
rect 337285 298696 337290 298752
rect 337346 298696 340124 298752
rect 337285 298694 340124 298696
rect 337285 298691 337351 298694
rect 583520 298604 584960 298844
rect 337745 298074 337811 298077
rect 337745 298072 340124 298074
rect 337745 298016 337750 298072
rect 337806 298016 340124 298072
rect 337745 298014 340124 298016
rect 337745 298011 337811 298014
rect 482829 297666 482895 297669
rect 479964 297664 482895 297666
rect 479964 297608 482834 297664
rect 482890 297608 482895 297664
rect 479964 297606 482895 297608
rect 482829 297603 482895 297606
rect 337653 297394 337719 297397
rect 337653 297392 340124 297394
rect 337653 297336 337658 297392
rect 337714 297336 340124 297392
rect 337653 297334 340124 297336
rect 337653 297331 337719 297334
rect 19374 296924 19380 296988
rect 19444 296986 19450 296988
rect 19793 296986 19859 296989
rect 19444 296984 19859 296986
rect 19444 296928 19798 296984
rect 19854 296928 19859 296984
rect 19444 296926 19859 296928
rect 19444 296924 19450 296926
rect 19793 296923 19859 296926
rect 19374 296788 19380 296852
rect 19444 296850 19450 296852
rect 20662 296850 20668 296852
rect 19444 296790 20668 296850
rect 19444 296788 19450 296790
rect 20662 296788 20668 296790
rect 20732 296788 20738 296852
rect 336917 296850 336983 296853
rect 336917 296848 340124 296850
rect 336917 296792 336922 296848
rect 336978 296792 340124 296848
rect 336917 296790 340124 296792
rect 336917 296787 336983 296790
rect 19374 296652 19380 296716
rect 19444 296714 19450 296716
rect 19444 296654 20730 296714
rect 19444 296652 19450 296654
rect 19374 296516 19380 296580
rect 19444 296578 19450 296580
rect 19793 296578 19859 296581
rect 20670 296580 20730 296654
rect 19444 296576 19859 296578
rect 19444 296520 19798 296576
rect 19854 296520 19859 296576
rect 19444 296518 19859 296520
rect 19444 296516 19450 296518
rect 19793 296515 19859 296518
rect 20662 296516 20668 296580
rect 20732 296516 20738 296580
rect 337653 296170 337719 296173
rect 337653 296168 340124 296170
rect 337653 296112 337658 296168
rect 337714 296112 340124 296168
rect 337653 296110 340124 296112
rect 337653 296107 337719 296110
rect 337101 295490 337167 295493
rect 337101 295488 340124 295490
rect 337101 295432 337106 295488
rect 337162 295432 340124 295488
rect 337101 295430 340124 295432
rect 337101 295427 337167 295430
rect 336917 294946 336983 294949
rect 336917 294944 340124 294946
rect 336917 294888 336922 294944
rect 336978 294888 340124 294944
rect 336917 294886 340124 294888
rect 336917 294883 336983 294886
rect 337653 294266 337719 294269
rect 337653 294264 340124 294266
rect 337653 294208 337658 294264
rect 337714 294208 340124 294264
rect 337653 294206 340124 294208
rect 337653 294203 337719 294206
rect 337653 293586 337719 293589
rect 337653 293584 340124 293586
rect 337653 293528 337658 293584
rect 337714 293528 340124 293584
rect 337653 293526 340124 293528
rect 337653 293523 337719 293526
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 482737 293042 482803 293045
rect 479964 293040 482803 293042
rect 479964 292984 482742 293040
rect 482798 292984 482803 293040
rect 479964 292982 482803 292984
rect 482737 292979 482803 292982
rect 337745 292906 337811 292909
rect 337745 292904 340124 292906
rect 337745 292848 337750 292904
rect 337806 292848 340124 292904
rect 337745 292846 340124 292848
rect 337745 292843 337811 292846
rect 337653 292362 337719 292365
rect 337653 292360 340124 292362
rect 337653 292304 337658 292360
rect 337714 292304 340124 292360
rect 337653 292302 340124 292304
rect 337653 292299 337719 292302
rect 337745 291682 337811 291685
rect 337745 291680 340124 291682
rect 337745 291624 337750 291680
rect 337806 291624 340124 291680
rect 337745 291622 340124 291624
rect 337745 291619 337811 291622
rect 48313 291138 48379 291141
rect 48630 291138 48636 291140
rect 48313 291136 48636 291138
rect 48313 291080 48318 291136
rect 48374 291080 48636 291136
rect 48313 291078 48636 291080
rect 48313 291075 48379 291078
rect 48630 291076 48636 291078
rect 48700 291076 48706 291140
rect 51022 291076 51028 291140
rect 51092 291138 51098 291140
rect 52361 291138 52427 291141
rect 51092 291136 52427 291138
rect 51092 291080 52366 291136
rect 52422 291080 52427 291136
rect 51092 291078 52427 291080
rect 51092 291076 51098 291078
rect 52361 291075 52427 291078
rect 53414 291076 53420 291140
rect 53484 291138 53490 291140
rect 53741 291138 53807 291141
rect 56501 291140 56567 291141
rect 56501 291138 56548 291140
rect 53484 291136 53807 291138
rect 53484 291080 53746 291136
rect 53802 291080 53807 291136
rect 53484 291078 53807 291080
rect 56456 291136 56548 291138
rect 56456 291080 56506 291136
rect 56456 291078 56548 291080
rect 53484 291076 53490 291078
rect 53741 291075 53807 291078
rect 56501 291076 56548 291078
rect 56612 291076 56618 291140
rect 58566 291076 58572 291140
rect 58636 291138 58642 291140
rect 59261 291138 59327 291141
rect 58636 291136 59327 291138
rect 58636 291080 59266 291136
rect 59322 291080 59327 291136
rect 58636 291078 59327 291080
rect 58636 291076 58642 291078
rect 56501 291075 56567 291076
rect 59261 291075 59327 291078
rect 61142 291076 61148 291140
rect 61212 291138 61218 291140
rect 62021 291138 62087 291141
rect 61212 291136 62087 291138
rect 61212 291080 62026 291136
rect 62082 291080 62087 291136
rect 61212 291078 62087 291080
rect 61212 291076 61218 291078
rect 62021 291075 62087 291078
rect 64086 291076 64092 291140
rect 64156 291138 64162 291140
rect 64781 291138 64847 291141
rect 64156 291136 64847 291138
rect 64156 291080 64786 291136
rect 64842 291080 64847 291136
rect 64156 291078 64847 291080
rect 64156 291076 64162 291078
rect 64781 291075 64847 291078
rect 68502 291076 68508 291140
rect 68572 291138 68578 291140
rect 68921 291138 68987 291141
rect 68572 291136 68987 291138
rect 68572 291080 68926 291136
rect 68982 291080 68987 291136
rect 68572 291078 68987 291080
rect 68572 291076 68578 291078
rect 68921 291075 68987 291078
rect 71078 291076 71084 291140
rect 71148 291138 71154 291140
rect 71681 291138 71747 291141
rect 71148 291136 71747 291138
rect 71148 291080 71686 291136
rect 71742 291080 71747 291136
rect 71148 291078 71747 291080
rect 71148 291076 71154 291078
rect 71681 291075 71747 291078
rect 76230 291076 76236 291140
rect 76300 291138 76306 291140
rect 77201 291138 77267 291141
rect 76300 291136 77267 291138
rect 76300 291080 77206 291136
rect 77262 291080 77267 291136
rect 76300 291078 77267 291080
rect 76300 291076 76306 291078
rect 77201 291075 77267 291078
rect 78438 291076 78444 291140
rect 78508 291138 78514 291140
rect 78581 291138 78647 291141
rect 78508 291136 78647 291138
rect 78508 291080 78586 291136
rect 78642 291080 78647 291136
rect 78508 291078 78647 291080
rect 78508 291076 78514 291078
rect 78581 291075 78647 291078
rect 81014 291076 81020 291140
rect 81084 291138 81090 291140
rect 81341 291138 81407 291141
rect 81084 291136 81407 291138
rect 81084 291080 81346 291136
rect 81402 291080 81407 291136
rect 81084 291078 81407 291080
rect 81084 291076 81090 291078
rect 81341 291075 81407 291078
rect 83590 291076 83596 291140
rect 83660 291138 83666 291140
rect 84101 291138 84167 291141
rect 83660 291136 84167 291138
rect 83660 291080 84106 291136
rect 84162 291080 84167 291136
rect 83660 291078 84167 291080
rect 83660 291076 83666 291078
rect 84101 291075 84167 291078
rect 86166 291076 86172 291140
rect 86236 291138 86242 291140
rect 86861 291138 86927 291141
rect 86236 291136 86927 291138
rect 86236 291080 86866 291136
rect 86922 291080 86927 291136
rect 86236 291078 86927 291080
rect 86236 291076 86242 291078
rect 86861 291075 86927 291078
rect 88558 291076 88564 291140
rect 88628 291138 88634 291140
rect 89621 291138 89687 291141
rect 91001 291140 91067 291141
rect 88628 291136 89687 291138
rect 88628 291080 89626 291136
rect 89682 291080 89687 291136
rect 88628 291078 89687 291080
rect 88628 291076 88634 291078
rect 89621 291075 89687 291078
rect 90950 291076 90956 291140
rect 91020 291138 91067 291140
rect 91020 291136 91112 291138
rect 91062 291080 91112 291136
rect 91020 291078 91112 291080
rect 91020 291076 91067 291078
rect 93526 291076 93532 291140
rect 93596 291138 93602 291140
rect 93761 291138 93827 291141
rect 93596 291136 93827 291138
rect 93596 291080 93766 291136
rect 93822 291080 93827 291136
rect 93596 291078 93827 291080
rect 93596 291076 93602 291078
rect 91001 291075 91067 291076
rect 93761 291075 93827 291078
rect 98678 291076 98684 291140
rect 98748 291138 98754 291140
rect 99281 291138 99347 291141
rect 98748 291136 99347 291138
rect 98748 291080 99286 291136
rect 99342 291080 99347 291136
rect 98748 291078 99347 291080
rect 98748 291076 98754 291078
rect 99281 291075 99347 291078
rect 106038 291076 106044 291140
rect 106108 291138 106114 291140
rect 106181 291138 106247 291141
rect 106108 291136 106247 291138
rect 106108 291080 106186 291136
rect 106242 291080 106247 291136
rect 106108 291078 106247 291080
rect 106108 291076 106114 291078
rect 106181 291075 106247 291078
rect 115974 291076 115980 291140
rect 116044 291138 116050 291140
rect 117221 291138 117287 291141
rect 116044 291136 117287 291138
rect 116044 291080 117226 291136
rect 117282 291080 117287 291136
rect 116044 291078 117287 291080
rect 116044 291076 116050 291078
rect 117221 291075 117287 291078
rect 208710 291076 208716 291140
rect 208780 291138 208786 291140
rect 209313 291138 209379 291141
rect 208780 291136 209379 291138
rect 208780 291080 209318 291136
rect 209374 291080 209379 291136
rect 208780 291078 209379 291080
rect 208780 291076 208786 291078
rect 209313 291075 209379 291078
rect 210734 291076 210740 291140
rect 210804 291138 210810 291140
rect 211061 291138 211127 291141
rect 210804 291136 211127 291138
rect 210804 291080 211066 291136
rect 211122 291080 211127 291136
rect 210804 291078 211127 291080
rect 210804 291076 210810 291078
rect 211061 291075 211127 291078
rect 213494 291076 213500 291140
rect 213564 291138 213570 291140
rect 213821 291138 213887 291141
rect 213564 291136 213887 291138
rect 213564 291080 213826 291136
rect 213882 291080 213887 291136
rect 213564 291078 213887 291080
rect 213564 291076 213570 291078
rect 213821 291075 213887 291078
rect 216254 291076 216260 291140
rect 216324 291138 216330 291140
rect 216489 291138 216555 291141
rect 216324 291136 216555 291138
rect 216324 291080 216494 291136
rect 216550 291080 216555 291136
rect 216324 291078 216555 291080
rect 216324 291076 216330 291078
rect 216489 291075 216555 291078
rect 218646 291076 218652 291140
rect 218716 291138 218722 291140
rect 219341 291138 219407 291141
rect 218716 291136 219407 291138
rect 218716 291080 219346 291136
rect 219402 291080 219407 291136
rect 218716 291078 219407 291080
rect 218716 291076 218722 291078
rect 219341 291075 219407 291078
rect 221038 291076 221044 291140
rect 221108 291138 221114 291140
rect 222101 291138 222167 291141
rect 223481 291140 223547 291141
rect 226241 291140 226307 291141
rect 221108 291136 222167 291138
rect 221108 291080 222106 291136
rect 222162 291080 222167 291136
rect 221108 291078 222167 291080
rect 221108 291076 221114 291078
rect 222101 291075 222167 291078
rect 223430 291076 223436 291140
rect 223500 291138 223547 291140
rect 223500 291136 223592 291138
rect 223542 291080 223592 291136
rect 223500 291078 223592 291080
rect 223500 291076 223547 291078
rect 226190 291076 226196 291140
rect 226260 291138 226307 291140
rect 226260 291136 226352 291138
rect 226302 291080 226352 291136
rect 226260 291078 226352 291080
rect 226260 291076 226307 291078
rect 228582 291076 228588 291140
rect 228652 291138 228658 291140
rect 228909 291138 228975 291141
rect 228652 291136 228975 291138
rect 228652 291080 228914 291136
rect 228970 291080 228975 291136
rect 228652 291078 228975 291080
rect 228652 291076 228658 291078
rect 223481 291075 223547 291076
rect 226241 291075 226307 291076
rect 228909 291075 228975 291078
rect 231158 291076 231164 291140
rect 231228 291138 231234 291140
rect 231761 291138 231827 291141
rect 231228 291136 231827 291138
rect 231228 291080 231766 291136
rect 231822 291080 231827 291136
rect 231228 291078 231827 291080
rect 231228 291076 231234 291078
rect 231761 291075 231827 291078
rect 238518 291076 238524 291140
rect 238588 291138 238594 291140
rect 238661 291138 238727 291141
rect 238588 291136 238727 291138
rect 238588 291080 238666 291136
rect 238722 291080 238727 291136
rect 238588 291078 238727 291080
rect 238588 291076 238594 291078
rect 238661 291075 238727 291078
rect 240910 291076 240916 291140
rect 240980 291138 240986 291140
rect 241421 291138 241487 291141
rect 240980 291136 241487 291138
rect 240980 291080 241426 291136
rect 241482 291080 241487 291136
rect 240980 291078 241487 291080
rect 240980 291076 240986 291078
rect 241421 291075 241487 291078
rect 244038 291076 244044 291140
rect 244108 291138 244114 291140
rect 244181 291138 244247 291141
rect 244108 291136 244247 291138
rect 244108 291080 244186 291136
rect 244242 291080 244247 291136
rect 244108 291078 244247 291080
rect 244108 291076 244114 291078
rect 244181 291075 244247 291078
rect 246062 291076 246068 291140
rect 246132 291138 246138 291140
rect 246941 291138 247007 291141
rect 246132 291136 247007 291138
rect 246132 291080 246946 291136
rect 247002 291080 247007 291136
rect 246132 291078 247007 291080
rect 246132 291076 246138 291078
rect 246941 291075 247007 291078
rect 248638 291076 248644 291140
rect 248708 291138 248714 291140
rect 249701 291138 249767 291141
rect 251081 291140 251147 291141
rect 248708 291136 249767 291138
rect 248708 291080 249706 291136
rect 249762 291080 249767 291136
rect 248708 291078 249767 291080
rect 248708 291076 248714 291078
rect 249701 291075 249767 291078
rect 251030 291076 251036 291140
rect 251100 291138 251147 291140
rect 251100 291136 251192 291138
rect 251142 291080 251192 291136
rect 251100 291078 251192 291080
rect 251100 291076 251147 291078
rect 253606 291076 253612 291140
rect 253676 291138 253682 291140
rect 253841 291138 253907 291141
rect 253676 291136 253907 291138
rect 253676 291080 253846 291136
rect 253902 291080 253907 291136
rect 253676 291078 253907 291080
rect 253676 291076 253682 291078
rect 251081 291075 251147 291076
rect 253841 291075 253907 291078
rect 255998 291076 256004 291140
rect 256068 291138 256074 291140
rect 256601 291138 256667 291141
rect 256068 291136 256667 291138
rect 256068 291080 256606 291136
rect 256662 291080 256667 291136
rect 256068 291078 256667 291080
rect 256068 291076 256074 291078
rect 256601 291075 256667 291078
rect 258574 291076 258580 291140
rect 258644 291138 258650 291140
rect 259361 291138 259427 291141
rect 258644 291136 259427 291138
rect 258644 291080 259366 291136
rect 259422 291080 259427 291136
rect 258644 291078 259427 291080
rect 258644 291076 258650 291078
rect 259361 291075 259427 291078
rect 263542 291076 263548 291140
rect 263612 291138 263618 291140
rect 264881 291138 264947 291141
rect 263612 291136 264947 291138
rect 263612 291080 264886 291136
rect 264942 291080 264947 291136
rect 263612 291078 264947 291080
rect 263612 291076 263618 291078
rect 264881 291075 264947 291078
rect 268510 291076 268516 291140
rect 268580 291138 268586 291140
rect 269021 291138 269087 291141
rect 268580 291136 269087 291138
rect 268580 291080 269026 291136
rect 269082 291080 269087 291136
rect 268580 291078 269087 291080
rect 268580 291076 268586 291078
rect 269021 291075 269087 291078
rect 271086 291076 271092 291140
rect 271156 291138 271162 291140
rect 271781 291138 271847 291141
rect 271156 291136 271847 291138
rect 271156 291080 271786 291136
rect 271842 291080 271847 291136
rect 271156 291078 271847 291080
rect 271156 291076 271162 291078
rect 271781 291075 271847 291078
rect 273662 291076 273668 291140
rect 273732 291138 273738 291140
rect 274541 291138 274607 291141
rect 273732 291136 274607 291138
rect 273732 291080 274546 291136
rect 274602 291080 274607 291136
rect 273732 291078 274607 291080
rect 273732 291076 273738 291078
rect 274541 291075 274607 291078
rect 276238 291076 276244 291140
rect 276308 291138 276314 291140
rect 277301 291138 277367 291141
rect 276308 291136 277367 291138
rect 276308 291080 277306 291136
rect 277362 291080 277367 291136
rect 276308 291078 277367 291080
rect 276308 291076 276314 291078
rect 277301 291075 277367 291078
rect 281022 291076 281028 291140
rect 281092 291138 281098 291140
rect 281441 291138 281507 291141
rect 281092 291136 281507 291138
rect 281092 291080 281446 291136
rect 281502 291080 281507 291136
rect 281092 291078 281507 291080
rect 281092 291076 281098 291078
rect 281441 291075 281507 291078
rect 283782 291076 283788 291140
rect 283852 291138 283858 291140
rect 284201 291138 284267 291141
rect 283852 291136 284267 291138
rect 283852 291080 284206 291136
rect 284262 291080 284267 291136
rect 283852 291078 284267 291080
rect 283852 291076 283858 291078
rect 284201 291075 284267 291078
rect 101070 290940 101076 291004
rect 101140 291002 101146 291004
rect 102041 291002 102107 291005
rect 101140 291000 102107 291002
rect 101140 290944 102046 291000
rect 102102 290944 102107 291000
rect 101140 290942 102107 290944
rect 101140 290940 101146 290942
rect 102041 290939 102107 290942
rect 113214 290940 113220 291004
rect 113284 291002 113290 291004
rect 114461 291002 114527 291005
rect 113284 291000 114527 291002
rect 113284 290944 114466 291000
rect 114522 290944 114527 291000
rect 113284 290942 114527 290944
rect 113284 290940 113290 290942
rect 114461 290939 114527 290942
rect 236494 290940 236500 291004
rect 236564 291002 236570 291004
rect 237281 291002 237347 291005
rect 236564 291000 237347 291002
rect 236564 290944 237286 291000
rect 237342 290944 237347 291000
rect 236564 290942 237347 290944
rect 236564 290940 236570 290942
rect 237281 290939 237347 290942
rect 337469 291002 337535 291005
rect 337469 291000 340124 291002
rect 337469 290944 337474 291000
rect 337530 290944 340124 291000
rect 337469 290942 340124 290944
rect 337469 290939 337535 290942
rect 111006 290804 111012 290868
rect 111076 290866 111082 290868
rect 111701 290866 111767 290869
rect 111076 290864 111767 290866
rect 111076 290808 111706 290864
rect 111762 290808 111767 290864
rect 111076 290806 111767 290808
rect 111076 290804 111082 290806
rect 111701 290803 111767 290806
rect 139710 290804 139716 290868
rect 139780 290866 139786 290868
rect 140681 290866 140747 290869
rect 139780 290864 140747 290866
rect 139780 290808 140686 290864
rect 140742 290808 140747 290864
rect 139780 290806 140747 290808
rect 139780 290804 139786 290806
rect 140681 290803 140747 290806
rect 64822 290668 64828 290732
rect 64892 290730 64898 290732
rect 66161 290730 66227 290733
rect 64892 290728 66227 290730
rect 64892 290672 66166 290728
rect 66222 290672 66227 290728
rect 64892 290670 66227 290672
rect 64892 290668 64898 290670
rect 66161 290667 66227 290670
rect 103830 290668 103836 290732
rect 103900 290730 103906 290732
rect 104801 290730 104867 290733
rect 118601 290732 118667 290733
rect 103900 290728 104867 290730
rect 103900 290672 104806 290728
rect 104862 290672 104867 290728
rect 103900 290670 104867 290672
rect 103900 290668 103906 290670
rect 104801 290667 104867 290670
rect 118550 290668 118556 290732
rect 118620 290730 118667 290732
rect 118620 290728 118712 290730
rect 118662 290672 118712 290728
rect 118620 290670 118712 290672
rect 118620 290668 118667 290670
rect 265934 290668 265940 290732
rect 266004 290730 266010 290732
rect 266261 290730 266327 290733
rect 266004 290728 266327 290730
rect 266004 290672 266266 290728
rect 266322 290672 266327 290728
rect 266004 290670 266327 290672
rect 266004 290668 266010 290670
rect 118601 290667 118667 290668
rect 266261 290667 266327 290670
rect 277342 290668 277348 290732
rect 277412 290730 277418 290732
rect 278681 290730 278747 290733
rect 277412 290728 278747 290730
rect 277412 290672 278686 290728
rect 278742 290672 278747 290728
rect 277412 290670 278747 290672
rect 277412 290668 277418 290670
rect 278681 290667 278747 290670
rect 126094 290396 126100 290460
rect 126164 290458 126170 290460
rect 126881 290458 126947 290461
rect 126164 290456 126947 290458
rect 126164 290400 126886 290456
rect 126942 290400 126947 290456
rect 126164 290398 126947 290400
rect 126164 290396 126170 290398
rect 126881 290395 126947 290398
rect 138422 290396 138428 290460
rect 138492 290458 138498 290460
rect 139301 290458 139367 290461
rect 138492 290456 139367 290458
rect 138492 290400 139306 290456
rect 139362 290400 139367 290456
rect 138492 290398 139367 290400
rect 138492 290396 138498 290398
rect 139301 290395 139367 290398
rect 260966 290396 260972 290460
rect 261036 290458 261042 290460
rect 262121 290458 262187 290461
rect 261036 290456 262187 290458
rect 261036 290400 262126 290456
rect 262182 290400 262187 290456
rect 261036 290398 262187 290400
rect 261036 290396 261042 290398
rect 262121 290395 262187 290398
rect 337101 290458 337167 290461
rect 337101 290456 340124 290458
rect 337101 290400 337106 290456
rect 337162 290400 340124 290456
rect 337101 290398 340124 290400
rect 337101 290395 337167 290398
rect 73470 290260 73476 290324
rect 73540 290322 73546 290324
rect 73981 290322 74047 290325
rect 73540 290320 74047 290322
rect 73540 290264 73986 290320
rect 74042 290264 74047 290320
rect 73540 290262 74047 290264
rect 73540 290260 73546 290262
rect 73981 290259 74047 290262
rect 120758 290260 120764 290324
rect 120828 290322 120834 290324
rect 121361 290322 121427 290325
rect 120828 290320 121427 290322
rect 120828 290264 121366 290320
rect 121422 290264 121427 290320
rect 120828 290262 121427 290264
rect 120828 290260 120834 290262
rect 121361 290259 121427 290262
rect 96286 290124 96292 290188
rect 96356 290186 96362 290188
rect 96521 290186 96587 290189
rect 96356 290184 96587 290186
rect 96356 290128 96526 290184
rect 96582 290128 96587 290184
rect 96356 290126 96587 290128
rect 96356 290124 96362 290126
rect 96521 290123 96587 290126
rect 108430 289988 108436 290052
rect 108500 290050 108506 290052
rect 108941 290050 109007 290053
rect 122833 290052 122899 290053
rect 108500 290048 109007 290050
rect 108500 289992 108946 290048
rect 109002 289992 109007 290048
rect 108500 289990 109007 289992
rect 108500 289988 108506 289990
rect 108941 289987 109007 289990
rect 122782 289988 122788 290052
rect 122852 290050 122899 290052
rect 122852 290048 122944 290050
rect 122894 289992 122944 290048
rect 122852 289990 122944 289992
rect 122852 289988 122899 289990
rect 233550 289988 233556 290052
rect 233620 290050 233626 290052
rect 234521 290050 234587 290053
rect 233620 290048 234587 290050
rect 233620 289992 234526 290048
rect 234582 289992 234587 290048
rect 233620 289990 234587 289992
rect 233620 289988 233626 289990
rect 122833 289987 122899 289988
rect 234521 289987 234587 289990
rect 286174 289852 286180 289916
rect 286244 289914 286250 289916
rect 286593 289914 286659 289917
rect 286244 289912 286659 289914
rect 286244 289856 286598 289912
rect 286654 289856 286659 289912
rect 286244 289854 286659 289856
rect 286244 289852 286250 289854
rect 286593 289851 286659 289854
rect 298502 289852 298508 289916
rect 298572 289914 298578 289916
rect 299013 289914 299079 289917
rect 299657 289916 299723 289917
rect 299606 289914 299612 289916
rect 298572 289912 299079 289914
rect 298572 289856 299018 289912
rect 299074 289856 299079 289912
rect 298572 289854 299079 289856
rect 299566 289854 299612 289914
rect 299676 289912 299723 289916
rect 299718 289856 299723 289912
rect 298572 289852 298578 289854
rect 299013 289851 299079 289854
rect 299606 289852 299612 289854
rect 299676 289852 299723 289856
rect 299657 289851 299723 289852
rect 310789 289916 310855 289917
rect 310789 289912 310836 289916
rect 310900 289914 310906 289916
rect 310789 289856 310794 289912
rect 310789 289852 310836 289856
rect 310900 289854 310946 289914
rect 310900 289852 310906 289854
rect 310789 289851 310855 289852
rect 337653 289778 337719 289781
rect 337653 289776 340124 289778
rect 337653 289720 337658 289776
rect 337714 289720 340124 289776
rect 337653 289718 340124 289720
rect 337653 289715 337719 289718
rect 3509 289098 3575 289101
rect 324957 289098 325023 289101
rect 3509 289096 325023 289098
rect 3509 289040 3514 289096
rect 3570 289040 324962 289096
rect 325018 289040 325023 289096
rect 3509 289038 325023 289040
rect 3509 289035 3575 289038
rect 324957 289035 325023 289038
rect 337745 289098 337811 289101
rect 337745 289096 340124 289098
rect 337745 289040 337750 289096
rect 337806 289040 340124 289096
rect 337745 289038 340124 289040
rect 337745 289035 337811 289038
rect 19374 288900 19380 288964
rect 19444 288962 19450 288964
rect 19742 288962 19748 288964
rect 19444 288902 19748 288962
rect 19444 288900 19450 288902
rect 19742 288900 19748 288902
rect 19812 288900 19818 288964
rect 178350 288764 178356 288828
rect 178420 288826 178426 288828
rect 179270 288826 179276 288828
rect 178420 288766 179276 288826
rect 178420 288764 178426 288766
rect 179270 288764 179276 288766
rect 179340 288764 179346 288828
rect 19374 288492 19380 288556
rect 19444 288554 19450 288556
rect 20846 288554 20852 288556
rect 19444 288494 20852 288554
rect 19444 288492 19450 288494
rect 20846 288492 20852 288494
rect 20916 288492 20922 288556
rect 337653 288418 337719 288421
rect 337653 288416 340124 288418
rect 337653 288360 337658 288416
rect 337714 288360 340124 288416
rect 337653 288358 340124 288360
rect 337653 288355 337719 288358
rect 482645 288282 482711 288285
rect 479964 288280 482711 288282
rect 479964 288224 482650 288280
rect 482706 288224 482711 288280
rect 479964 288222 482711 288224
rect 482645 288219 482711 288222
rect 179270 287812 179276 287876
rect 179340 287874 179346 287876
rect 179638 287874 179644 287876
rect 179340 287814 179644 287874
rect 179340 287812 179346 287814
rect 179638 287812 179644 287814
rect 179708 287812 179714 287876
rect 337745 287874 337811 287877
rect 337745 287872 340124 287874
rect 337745 287816 337750 287872
rect 337806 287816 340124 287872
rect 337745 287814 340124 287816
rect 337745 287811 337811 287814
rect 18454 287676 18460 287740
rect 18524 287738 18530 287740
rect 46197 287738 46263 287741
rect 18524 287736 46263 287738
rect 18524 287680 46202 287736
rect 46258 287680 46263 287736
rect 18524 287678 46263 287680
rect 18524 287676 18530 287678
rect 46197 287675 46263 287678
rect 179638 287676 179644 287740
rect 179708 287738 179714 287740
rect 180006 287738 180012 287740
rect 179708 287678 180012 287738
rect 179708 287676 179714 287678
rect 180006 287676 180012 287678
rect 180076 287676 180082 287740
rect 150893 287468 150959 287469
rect 150832 287466 150838 287468
rect 150802 287406 150838 287466
rect 150902 287464 150959 287468
rect 150954 287408 150959 287464
rect 150832 287404 150838 287406
rect 150902 287404 150959 287408
rect 150893 287403 150959 287404
rect 180333 287466 180399 287469
rect 180558 287466 180564 287468
rect 180333 287464 180564 287466
rect 180333 287408 180338 287464
rect 180394 287408 180564 287464
rect 180333 287406 180564 287408
rect 180333 287403 180399 287406
rect 180558 287404 180564 287406
rect 180628 287404 180634 287468
rect 336917 287194 336983 287197
rect 336917 287192 340124 287194
rect 336917 287136 336922 287192
rect 336978 287136 340124 287192
rect 336917 287134 340124 287136
rect 336917 287131 336983 287134
rect 337469 286922 337535 286925
rect 337150 286920 337535 286922
rect 337150 286864 337474 286920
rect 337530 286864 337535 286920
rect 337150 286862 337535 286864
rect 337150 286789 337210 286862
rect 337469 286859 337535 286862
rect 337101 286784 337210 286789
rect 337101 286728 337106 286784
rect 337162 286728 337210 286784
rect 337101 286726 337210 286728
rect 337101 286723 337167 286726
rect 336733 286514 336799 286517
rect 336733 286512 340124 286514
rect 336733 286456 336738 286512
rect 336794 286456 340124 286512
rect 336733 286454 340124 286456
rect 336733 286451 336799 286454
rect 337469 285834 337535 285837
rect 337469 285832 340124 285834
rect 337469 285776 337474 285832
rect 337530 285776 340124 285832
rect 337469 285774 340124 285776
rect 337469 285771 337535 285774
rect 337285 285290 337351 285293
rect 337285 285288 340124 285290
rect 337285 285232 337290 285288
rect 337346 285232 340124 285288
rect 583520 285276 584960 285516
rect 337285 285230 340124 285232
rect 337285 285227 337351 285230
rect 337653 284610 337719 284613
rect 337653 284608 340124 284610
rect 337653 284552 337658 284608
rect 337714 284552 340124 284608
rect 337653 284550 340124 284552
rect 337653 284547 337719 284550
rect 337653 283930 337719 283933
rect 337653 283928 340124 283930
rect 337653 283872 337658 283928
rect 337714 283872 340124 283928
rect 337653 283870 340124 283872
rect 337653 283867 337719 283870
rect 482553 283658 482619 283661
rect 479964 283656 482619 283658
rect 479964 283600 482558 283656
rect 482614 283600 482619 283656
rect 479964 283598 482619 283600
rect 482553 283595 482619 283598
rect 337745 283386 337811 283389
rect 337745 283384 340124 283386
rect 337745 283328 337750 283384
rect 337806 283328 340124 283384
rect 337745 283326 340124 283328
rect 337745 283323 337811 283326
rect 160001 283250 160067 283253
rect 319437 283250 319503 283253
rect 157198 283248 160067 283250
rect 157198 283220 160006 283248
rect 156588 283192 160006 283220
rect 160062 283192 160067 283248
rect 317094 283248 319503 283250
rect 317094 283220 319442 283248
rect 156588 283190 160067 283192
rect 156588 283160 157258 283190
rect 160001 283187 160067 283190
rect 316572 283192 319442 283220
rect 319498 283192 319503 283248
rect 316572 283190 319503 283192
rect 316572 283160 317154 283190
rect 319437 283187 319503 283190
rect 337653 282706 337719 282709
rect 337653 282704 340124 282706
rect 337653 282648 337658 282704
rect 337714 282648 340124 282704
rect 337653 282646 340124 282648
rect 337653 282643 337719 282646
rect 337745 282026 337811 282029
rect 337745 282024 340124 282026
rect 337745 281968 337750 282024
rect 337806 281968 340124 282024
rect 337745 281966 340124 281968
rect 337745 281963 337811 281966
rect 337653 281346 337719 281349
rect 337653 281344 340124 281346
rect 337653 281288 337658 281344
rect 337714 281288 340124 281344
rect 337653 281286 340124 281288
rect 337653 281283 337719 281286
rect 336273 280802 336339 280805
rect 336273 280800 340124 280802
rect 336273 280744 336278 280800
rect 336334 280744 340124 280800
rect 336273 280742 340124 280744
rect 336273 280739 336339 280742
rect -960 279972 480 280212
rect 336825 280122 336891 280125
rect 336825 280120 340124 280122
rect 336825 280064 336830 280120
rect 336886 280064 340124 280120
rect 336825 280062 340124 280064
rect 336825 280059 336891 280062
rect 336733 279442 336799 279445
rect 336733 279440 340124 279442
rect 336733 279384 336738 279440
rect 336794 279384 340124 279440
rect 336733 279382 340124 279384
rect 336733 279379 336799 279382
rect 482461 279034 482527 279037
rect 479964 279032 482527 279034
rect 479964 278976 482466 279032
rect 482522 278976 482527 279032
rect 479964 278974 482527 278976
rect 482461 278971 482527 278974
rect 337745 278898 337811 278901
rect 337745 278896 340124 278898
rect 337745 278840 337750 278896
rect 337806 278840 340124 278896
rect 337745 278838 340124 278840
rect 337745 278835 337811 278838
rect 337653 278218 337719 278221
rect 337653 278216 340124 278218
rect 337653 278160 337658 278216
rect 337714 278160 340124 278216
rect 337653 278158 340124 278160
rect 337653 278155 337719 278158
rect 337009 277538 337075 277541
rect 337193 277538 337259 277541
rect 337009 277536 337259 277538
rect 337009 277480 337014 277536
rect 337070 277480 337198 277536
rect 337254 277480 337259 277536
rect 337009 277478 337259 277480
rect 337009 277475 337075 277478
rect 337193 277475 337259 277478
rect 337745 277538 337811 277541
rect 337745 277536 340124 277538
rect 337745 277480 337750 277536
rect 337806 277480 340124 277536
rect 337745 277478 340124 277480
rect 337745 277475 337811 277478
rect 337009 277402 337075 277405
rect 337285 277402 337351 277405
rect 337837 277402 337903 277405
rect 337009 277400 337351 277402
rect 337009 277344 337014 277400
rect 337070 277344 337290 277400
rect 337346 277344 337351 277400
rect 337009 277342 337351 277344
rect 337009 277339 337075 277342
rect 337285 277339 337351 277342
rect 337702 277400 337903 277402
rect 337702 277344 337842 277400
rect 337898 277344 337903 277400
rect 337702 277342 337903 277344
rect 337285 277266 337351 277269
rect 337702 277266 337762 277342
rect 337837 277339 337903 277342
rect 337285 277264 337762 277266
rect 337285 277208 337290 277264
rect 337346 277208 337762 277264
rect 337285 277206 337762 277208
rect 337285 277203 337351 277206
rect 337837 276858 337903 276861
rect 337837 276856 340124 276858
rect 337837 276800 337842 276856
rect 337898 276800 340124 276856
rect 337837 276798 340124 276800
rect 337837 276795 337903 276798
rect 337377 276314 337443 276317
rect 337377 276312 340124 276314
rect 337377 276256 337382 276312
rect 337438 276256 340124 276312
rect 337377 276254 340124 276256
rect 337377 276251 337443 276254
rect 337837 275634 337903 275637
rect 337837 275632 340124 275634
rect 337837 275576 337842 275632
rect 337898 275576 340124 275632
rect 337837 275574 340124 275576
rect 337837 275571 337903 275574
rect 337377 274954 337443 274957
rect 337377 274952 340124 274954
rect 337377 274896 337382 274952
rect 337438 274896 340124 274952
rect 337377 274894 340124 274896
rect 337377 274891 337443 274894
rect 337101 274410 337167 274413
rect 337101 274408 340124 274410
rect 337101 274352 337106 274408
rect 337162 274352 340124 274408
rect 337101 274350 340124 274352
rect 337101 274347 337167 274350
rect 482369 274274 482435 274277
rect 479964 274272 482435 274274
rect 479964 274216 482374 274272
rect 482430 274216 482435 274272
rect 479964 274214 482435 274216
rect 482369 274211 482435 274214
rect 337837 273730 337903 273733
rect 337837 273728 340124 273730
rect 337837 273672 337842 273728
rect 337898 273672 340124 273728
rect 337837 273670 340124 273672
rect 337837 273667 337903 273670
rect 337193 273050 337259 273053
rect 337193 273048 340124 273050
rect 337193 272992 337198 273048
rect 337254 272992 340124 273048
rect 337193 272990 340124 272992
rect 337193 272987 337259 272990
rect 337837 272370 337903 272373
rect 337837 272368 340124 272370
rect 337837 272312 337842 272368
rect 337898 272312 340124 272368
rect 337837 272310 340124 272312
rect 337837 272307 337903 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 337101 271826 337167 271829
rect 337101 271824 340124 271826
rect 337101 271768 337106 271824
rect 337162 271768 340124 271824
rect 337101 271766 340124 271768
rect 337101 271763 337167 271766
rect 337837 271146 337903 271149
rect 337837 271144 340124 271146
rect 337837 271088 337842 271144
rect 337898 271088 340124 271144
rect 337837 271086 340124 271088
rect 337837 271083 337903 271086
rect 336181 270466 336247 270469
rect 336181 270464 340124 270466
rect 336181 270408 336186 270464
rect 336242 270408 340124 270464
rect 336181 270406 340124 270408
rect 336181 270403 336247 270406
rect 337837 269786 337903 269789
rect 337837 269784 340124 269786
rect 337837 269728 337842 269784
rect 337898 269728 340124 269784
rect 337837 269726 340124 269728
rect 337837 269723 337903 269726
rect 482369 269650 482435 269653
rect 479964 269648 482435 269650
rect 479964 269592 482374 269648
rect 482430 269592 482435 269648
rect 479964 269590 482435 269592
rect 482369 269587 482435 269590
rect 337009 269242 337075 269245
rect 337009 269240 340124 269242
rect 337009 269184 337014 269240
rect 337070 269184 340124 269240
rect 337009 269182 340124 269184
rect 337009 269179 337075 269182
rect 337285 268562 337351 268565
rect 337285 268560 340124 268562
rect 337285 268504 337290 268560
rect 337346 268504 340124 268560
rect 337285 268502 340124 268504
rect 337285 268499 337351 268502
rect 338021 267882 338087 267885
rect 338021 267880 340124 267882
rect 338021 267824 338026 267880
rect 338082 267824 340124 267880
rect 338021 267822 340124 267824
rect 338021 267819 338087 267822
rect 178166 267684 178172 267748
rect 178236 267746 178242 267748
rect 178677 267746 178743 267749
rect 178236 267744 178743 267746
rect 178236 267688 178682 267744
rect 178738 267688 178743 267744
rect 178236 267686 178743 267688
rect 178236 267684 178242 267686
rect 178677 267683 178743 267686
rect 337929 267338 337995 267341
rect 337929 267336 340124 267338
rect -960 267052 480 267292
rect 337929 267280 337934 267336
rect 337990 267280 340124 267336
rect 337929 267278 340124 267280
rect 337929 267275 337995 267278
rect 337745 266658 337811 266661
rect 337745 266656 340124 266658
rect 337745 266600 337750 266656
rect 337806 266600 340124 266656
rect 337745 266598 340124 266600
rect 337745 266595 337811 266598
rect 337653 265978 337719 265981
rect 337653 265976 340124 265978
rect 337653 265920 337658 265976
rect 337714 265920 340124 265976
rect 337653 265918 340124 265920
rect 337653 265915 337719 265918
rect 337469 265298 337535 265301
rect 337469 265296 340124 265298
rect 337469 265240 337474 265296
rect 337530 265240 340124 265296
rect 337469 265238 340124 265240
rect 337469 265235 337535 265238
rect 481909 265026 481975 265029
rect 479964 265024 481975 265026
rect 479964 264968 481914 265024
rect 481970 264968 481975 265024
rect 479964 264966 481975 264968
rect 481909 264963 481975 264966
rect 337561 264754 337627 264757
rect 337561 264752 340124 264754
rect 337561 264696 337566 264752
rect 337622 264696 340124 264752
rect 337561 264694 340124 264696
rect 337561 264691 337627 264694
rect 336825 264074 336891 264077
rect 336825 264072 340124 264074
rect 336825 264016 336830 264072
rect 336886 264016 340124 264072
rect 336825 264014 340124 264016
rect 336825 264011 336891 264014
rect 337469 263394 337535 263397
rect 337469 263392 340124 263394
rect 337469 263336 337474 263392
rect 337530 263336 340124 263392
rect 337469 263334 340124 263336
rect 337469 263331 337535 263334
rect 337377 262850 337443 262853
rect 337377 262848 340124 262850
rect 337377 262792 337382 262848
rect 337438 262792 340124 262848
rect 337377 262790 340124 262792
rect 337377 262787 337443 262790
rect 337469 262170 337535 262173
rect 337469 262168 340124 262170
rect 337469 262112 337474 262168
rect 337530 262112 340124 262168
rect 337469 262110 340124 262112
rect 337469 262107 337535 262110
rect 337653 261490 337719 261493
rect 337653 261488 340124 261490
rect 337653 261432 337658 261488
rect 337714 261432 340124 261488
rect 337653 261430 340124 261432
rect 337653 261427 337719 261430
rect 337745 260810 337811 260813
rect 337745 260808 340124 260810
rect 337745 260752 337750 260808
rect 337806 260752 340124 260808
rect 337745 260750 340124 260752
rect 337745 260747 337811 260750
rect 482277 260402 482343 260405
rect 479964 260400 482343 260402
rect 479964 260344 482282 260400
rect 482338 260344 482343 260400
rect 479964 260342 482343 260344
rect 482277 260339 482343 260342
rect 337653 260266 337719 260269
rect 337653 260264 340124 260266
rect 337653 260208 337658 260264
rect 337714 260208 340124 260264
rect 337653 260206 340124 260208
rect 337653 260203 337719 260206
rect 337101 259586 337167 259589
rect 337101 259584 340124 259586
rect 337101 259528 337106 259584
rect 337162 259528 340124 259584
rect 337101 259526 340124 259528
rect 337101 259523 337167 259526
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 339033 258634 339099 258637
rect 340094 258634 340154 258876
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 339033 258632 340154 258634
rect 339033 258576 339038 258632
rect 339094 258576 340154 258632
rect 339033 258574 340154 258576
rect 339033 258571 339099 258574
rect 337653 258362 337719 258365
rect 337653 258360 340124 258362
rect 337653 258304 337658 258360
rect 337714 258304 340124 258360
rect 337653 258302 340124 258304
rect 337653 258299 337719 258302
rect 178166 258164 178172 258228
rect 178236 258226 178242 258228
rect 178236 258166 178602 258226
rect 178236 258164 178242 258166
rect 178166 257892 178172 257956
rect 178236 257954 178242 257956
rect 178542 257954 178602 258166
rect 178236 257894 178602 257954
rect 178236 257892 178242 257894
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 177389 253874 177455 253877
rect 178166 253874 178172 253876
rect 177389 253872 178172 253874
rect 177389 253816 177394 253872
rect 177450 253816 178172 253872
rect 177389 253814 178172 253816
rect 177389 253811 177455 253814
rect 178166 253812 178172 253814
rect 178236 253812 178242 253876
rect 179822 245924 179828 245988
rect 179892 245924 179898 245988
rect 179830 245716 179890 245924
rect 179822 245652 179828 245716
rect 179892 245652 179898 245716
rect 583520 245428 584960 245668
rect 179638 244700 179644 244764
rect 179708 244762 179714 244764
rect 179708 244702 179890 244762
rect 179708 244700 179714 244702
rect 179270 244564 179276 244628
rect 179340 244626 179346 244628
rect 179340 244566 179706 244626
rect 179340 244564 179346 244566
rect 179646 244356 179706 244566
rect 177757 244290 177823 244293
rect 178350 244292 178356 244356
rect 178420 244354 178426 244356
rect 179270 244354 179276 244356
rect 178420 244294 179276 244354
rect 178420 244292 178426 244294
rect 179270 244292 179276 244294
rect 179340 244292 179346 244356
rect 179638 244292 179644 244356
rect 179708 244292 179714 244356
rect 177622 244288 177823 244290
rect 177622 244232 177762 244288
rect 177818 244232 177823 244288
rect 177622 244230 177823 244232
rect 177389 244082 177455 244085
rect 177622 244082 177682 244230
rect 177757 244227 177823 244230
rect 179830 244218 179890 244702
rect 177389 244080 177682 244082
rect 177389 244024 177394 244080
rect 177450 244024 177682 244080
rect 177389 244022 177682 244024
rect 179278 244158 179890 244218
rect 177389 244019 177455 244022
rect 179278 243810 179338 244158
rect 179597 243948 179663 243949
rect 179597 243946 179644 243948
rect 179552 243944 179644 243946
rect 179552 243888 179602 243944
rect 179552 243886 179644 243888
rect 179597 243884 179644 243886
rect 179708 243884 179714 243948
rect 179822 243884 179828 243948
rect 179892 243884 179898 243948
rect 179597 243883 179663 243884
rect 179638 243810 179644 243812
rect 179278 243750 179644 243810
rect 179638 243748 179644 243750
rect 179708 243748 179714 243812
rect 179830 243676 179890 243884
rect 179822 243612 179828 243676
rect 179892 243612 179898 243676
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 16849 240954 16915 240957
rect 177205 240954 177271 240957
rect 16849 240952 19442 240954
rect 16849 240896 16854 240952
rect 16910 240924 19442 240952
rect 177205 240952 179522 240954
rect 16910 240896 20056 240924
rect 16849 240894 20056 240896
rect 16849 240891 16915 240894
rect 19382 240864 20056 240894
rect 177205 240896 177210 240952
rect 177266 240924 179522 240952
rect 177266 240896 180032 240924
rect 177205 240894 180032 240896
rect 177205 240891 177271 240894
rect 179462 240864 180032 240894
rect 16757 240002 16823 240005
rect 177297 240002 177363 240005
rect 16757 240000 19442 240002
rect 16757 239944 16762 240000
rect 16818 239972 19442 240000
rect 177297 240000 179522 240002
rect 16818 239944 20056 239972
rect 16757 239942 20056 239944
rect 16757 239939 16823 239942
rect 19382 239912 20056 239942
rect 177297 239944 177302 240000
rect 177358 239972 179522 240000
rect 177358 239944 180032 239972
rect 177297 239942 180032 239944
rect 177297 239939 177363 239942
rect 179462 239912 180032 239942
rect 178350 239396 178356 239460
rect 178420 239458 178426 239460
rect 179270 239458 179276 239460
rect 178420 239398 179276 239458
rect 178420 239396 178426 239398
rect 179270 239396 179276 239398
rect 179340 239396 179346 239460
rect 17769 237826 17835 237829
rect 177389 237826 177455 237829
rect 17769 237824 19442 237826
rect 17769 237768 17774 237824
rect 17830 237796 19442 237824
rect 177389 237824 179522 237826
rect 17830 237768 20056 237796
rect 17769 237766 20056 237768
rect 17769 237763 17835 237766
rect 19382 237736 20056 237766
rect 177389 237768 177394 237824
rect 177450 237796 179522 237824
rect 177450 237768 180032 237796
rect 177389 237766 180032 237768
rect 177389 237763 177455 237766
rect 179462 237736 180032 237766
rect 17677 236874 17743 236877
rect 177481 236874 177547 236877
rect 17677 236872 19442 236874
rect 17677 236816 17682 236872
rect 17738 236844 19442 236872
rect 177481 236872 179522 236874
rect 17738 236816 20056 236844
rect 17677 236814 20056 236816
rect 17677 236811 17743 236814
rect 19382 236784 20056 236814
rect 177481 236816 177486 236872
rect 177542 236844 179522 236872
rect 177542 236816 180032 236844
rect 177481 236814 180032 236816
rect 177481 236811 177547 236814
rect 179462 236784 180032 236814
rect 179270 236540 179276 236604
rect 179340 236602 179346 236604
rect 179638 236602 179644 236604
rect 179340 236542 179644 236602
rect 179340 236540 179346 236542
rect 179638 236540 179644 236542
rect 179708 236540 179714 236604
rect 179597 236468 179663 236469
rect 179597 236466 179644 236468
rect 179552 236464 179644 236466
rect 179552 236408 179602 236464
rect 179552 236406 179644 236408
rect 179597 236404 179644 236406
rect 179708 236404 179714 236468
rect 179597 236403 179663 236404
rect 17493 235106 17559 235109
rect 177665 235106 177731 235109
rect 17493 235104 19442 235106
rect 17493 235048 17498 235104
rect 17554 235076 19442 235104
rect 177665 235104 179522 235106
rect 17554 235048 20056 235076
rect 17493 235046 20056 235048
rect 17493 235043 17559 235046
rect 19382 235016 20056 235046
rect 177665 235048 177670 235104
rect 177726 235076 179522 235104
rect 177726 235048 180032 235076
rect 177665 235046 180032 235048
rect 177665 235043 177731 235046
rect 179462 235016 180032 235046
rect 179270 234772 179276 234836
rect 179340 234834 179346 234836
rect 179340 234774 179522 234834
rect 179340 234772 179346 234774
rect 177757 234698 177823 234701
rect 179270 234698 179276 234700
rect 177757 234696 179276 234698
rect 177757 234640 177762 234696
rect 177818 234640 179276 234696
rect 177757 234638 179276 234640
rect 177757 234635 177823 234638
rect 179270 234636 179276 234638
rect 179340 234636 179346 234700
rect 178166 234364 178172 234428
rect 178236 234426 178242 234428
rect 179270 234426 179276 234428
rect 178236 234366 179276 234426
rect 178236 234364 178242 234366
rect 179270 234364 179276 234366
rect 179340 234364 179346 234428
rect 179270 234228 179276 234292
rect 179340 234290 179346 234292
rect 179462 234290 179522 234774
rect 179340 234230 179522 234290
rect 179340 234228 179346 234230
rect 17401 234018 17467 234021
rect 177573 234018 177639 234021
rect 17401 234016 19442 234018
rect 17401 233960 17406 234016
rect 17462 233988 19442 234016
rect 177573 234016 179522 234018
rect 17462 233960 20056 233988
rect 17401 233958 20056 233960
rect 17401 233955 17467 233958
rect 19382 233928 20056 233958
rect 177573 233960 177578 234016
rect 177634 233988 179522 234016
rect 177634 233960 180032 233988
rect 177573 233958 180032 233960
rect 177573 233955 177639 233958
rect 179462 233928 180032 233958
rect 179454 233004 179460 233068
rect 179524 233004 179530 233068
rect 179638 233004 179644 233068
rect 179708 233004 179714 233068
rect 179822 233004 179828 233068
rect 179892 233004 179898 233068
rect 179462 232796 179522 233004
rect 179646 232796 179706 233004
rect 179830 232796 179890 233004
rect 179454 232732 179460 232796
rect 179524 232732 179530 232796
rect 179638 232732 179644 232796
rect 179708 232732 179714 232796
rect 179822 232732 179828 232796
rect 179892 232732 179898 232796
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 17585 232250 17651 232253
rect 177113 232250 177179 232253
rect 177757 232250 177823 232253
rect 17585 232248 19442 232250
rect 17585 232192 17590 232248
rect 17646 232220 19442 232248
rect 177113 232248 179522 232250
rect 17646 232192 20056 232220
rect 17585 232190 20056 232192
rect 17585 232187 17651 232190
rect 19382 232160 20056 232190
rect 177113 232192 177118 232248
rect 177174 232192 177762 232248
rect 177818 232220 179522 232248
rect 583520 232236 584960 232326
rect 177818 232192 180032 232220
rect 177113 232190 180032 232192
rect 177113 232187 177179 232190
rect 177757 232187 177823 232190
rect 179462 232160 180032 232190
rect -960 227884 480 228124
rect 178166 224844 178172 224908
rect 178236 224906 178242 224908
rect 179454 224906 179460 224908
rect 178236 224846 179460 224906
rect 178236 224844 178242 224846
rect 179454 224844 179460 224846
rect 179524 224844 179530 224908
rect 179638 224844 179644 224908
rect 179708 224844 179714 224908
rect 177982 224708 177988 224772
rect 178052 224770 178058 224772
rect 179454 224770 179460 224772
rect 178052 224710 179460 224770
rect 178052 224708 178058 224710
rect 179454 224708 179460 224710
rect 179524 224708 179530 224772
rect 179646 224636 179706 224844
rect 179638 224572 179644 224636
rect 179708 224572 179714 224636
rect 159081 223410 159147 223413
rect 159357 223410 159423 223413
rect 317413 223410 317479 223413
rect 319897 223410 319963 223413
rect 157198 223408 159423 223410
rect 157198 223380 159086 223408
rect 156588 223352 159086 223380
rect 159142 223352 159362 223408
rect 159418 223352 159423 223408
rect 317094 223408 319963 223410
rect 317094 223380 317418 223408
rect 156588 223350 159423 223352
rect 156588 223320 157258 223350
rect 159081 223347 159147 223350
rect 159357 223347 159423 223350
rect 316572 223352 317418 223380
rect 317474 223352 319902 223408
rect 319958 223352 319963 223408
rect 316572 223350 319963 223352
rect 316572 223320 317154 223350
rect 317413 223347 317479 223350
rect 319897 223347 319963 223350
rect 177798 222668 177804 222732
rect 177868 222730 177874 222732
rect 179270 222730 179276 222732
rect 177868 222670 179276 222730
rect 177868 222668 177874 222670
rect 179270 222668 179276 222670
rect 179340 222668 179346 222732
rect 158713 221778 158779 221781
rect 159449 221778 159515 221781
rect 317505 221778 317571 221781
rect 319621 221778 319687 221781
rect 157198 221776 159515 221778
rect 157198 221748 158718 221776
rect 156588 221720 158718 221748
rect 158774 221720 159454 221776
rect 159510 221720 159515 221776
rect 317094 221776 319687 221778
rect 317094 221748 317510 221776
rect 156588 221718 159515 221720
rect 156588 221688 157258 221718
rect 158713 221715 158779 221718
rect 159449 221715 159515 221718
rect 316572 221720 317510 221748
rect 317566 221720 319626 221776
rect 319682 221720 319687 221776
rect 316572 221718 319687 221720
rect 316572 221688 317154 221718
rect 317505 221715 317571 221718
rect 319621 221715 319687 221718
rect 318793 220826 318859 220829
rect 319713 220826 319779 220829
rect 318793 220824 319779 220826
rect 318793 220768 318798 220824
rect 318854 220768 319718 220824
rect 319774 220768 319779 220824
rect 318793 220766 319779 220768
rect 318793 220763 318859 220766
rect 319713 220763 319779 220766
rect 158805 220418 158871 220421
rect 318793 220418 318859 220421
rect 157198 220416 158871 220418
rect 157198 220388 158810 220416
rect 156588 220360 158810 220388
rect 158866 220360 158871 220416
rect 317094 220416 318859 220418
rect 317094 220388 318798 220416
rect 156588 220358 158871 220360
rect 156588 220328 157258 220358
rect 158805 220355 158871 220358
rect 316572 220360 318798 220388
rect 318854 220360 318859 220416
rect 316572 220358 318859 220360
rect 316572 220328 317154 220358
rect 318793 220355 318859 220358
rect 178350 220084 178356 220148
rect 178420 220146 178426 220148
rect 179270 220146 179276 220148
rect 178420 220086 179276 220146
rect 178420 220084 178426 220086
rect 179270 220084 179276 220086
rect 179340 220084 179346 220148
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 158989 218922 159055 218925
rect 318885 218922 318951 218925
rect 157198 218920 159055 218922
rect 157198 218892 158994 218920
rect 156588 218864 158994 218892
rect 159050 218864 159055 218920
rect 317094 218920 318951 218922
rect 317094 218892 318890 218920
rect 156588 218862 159055 218864
rect 156588 218832 157258 218862
rect 158989 218859 159055 218862
rect 316572 218864 318890 218892
rect 318946 218864 318951 218920
rect 583520 218908 584960 218998
rect 316572 218862 318951 218864
rect 316572 218832 317154 218862
rect 318885 218859 318951 218862
rect 318885 218106 318951 218109
rect 319805 218106 319871 218109
rect 318885 218104 319871 218106
rect 318885 218048 318890 218104
rect 318946 218048 319810 218104
rect 319866 218048 319871 218104
rect 318885 218046 319871 218048
rect 318885 218043 318951 218046
rect 319805 218043 319871 218046
rect 158897 217698 158963 217701
rect 317597 217698 317663 217701
rect 319437 217698 319503 217701
rect 157198 217696 158963 217698
rect 157198 217668 158902 217696
rect 156588 217640 158902 217668
rect 158958 217640 158963 217696
rect 317094 217696 319503 217698
rect 317094 217668 317602 217696
rect 156588 217638 158963 217640
rect 156588 217608 157258 217638
rect 158897 217635 158963 217638
rect 316572 217640 317602 217668
rect 317658 217640 319442 217696
rect 319498 217640 319503 217696
rect 316572 217638 319503 217640
rect 316572 217608 317154 217638
rect 317597 217635 317663 217638
rect 319437 217635 319503 217638
rect 158897 216746 158963 216749
rect 159541 216746 159607 216749
rect 158897 216744 159607 216746
rect 158897 216688 158902 216744
rect 158958 216688 159546 216744
rect 159602 216688 159607 216744
rect 158897 216686 159607 216688
rect 158897 216683 158963 216686
rect 159541 216683 159607 216686
rect -960 214828 480 215068
rect 16941 214026 17007 214029
rect 177849 214026 177915 214029
rect 16941 214024 19442 214026
rect 16941 213968 16946 214024
rect 17002 213996 19442 214024
rect 177849 214024 179522 214026
rect 17002 213968 20056 213996
rect 16941 213966 20056 213968
rect 16941 213963 17007 213966
rect 19382 213936 20056 213966
rect 177849 213968 177854 214024
rect 177910 213996 179522 214024
rect 177910 213968 180032 213996
rect 177849 213966 180032 213968
rect 177849 213963 177915 213966
rect 179462 213936 180032 213966
rect 17861 212394 17927 212397
rect 177021 212394 177087 212397
rect 17861 212392 19442 212394
rect 17861 212336 17866 212392
rect 17922 212364 19442 212392
rect 177021 212392 179522 212394
rect 17922 212336 20056 212364
rect 17861 212334 20056 212336
rect 17861 212331 17927 212334
rect 19382 212304 20056 212334
rect 177021 212336 177026 212392
rect 177082 212364 179522 212392
rect 177082 212336 180032 212364
rect 177021 212334 180032 212336
rect 177021 212331 177087 212334
rect 179462 212304 180032 212334
rect 16941 212122 17007 212125
rect 177849 212122 177915 212125
rect 16941 212120 19442 212122
rect 16941 212064 16946 212120
rect 17002 212092 19442 212120
rect 177849 212120 179522 212122
rect 17002 212064 20056 212092
rect 16941 212062 20056 212064
rect 16941 212059 17007 212062
rect 19382 212032 20056 212062
rect 177849 212064 177854 212120
rect 177910 212092 179522 212120
rect 177910 212064 180032 212092
rect 177849 212062 180032 212064
rect 177849 212059 177915 212062
rect 179462 212032 180032 212062
rect 179822 210564 179828 210628
rect 179892 210564 179898 210628
rect 179638 210292 179644 210356
rect 179708 210354 179714 210356
rect 179830 210354 179890 210564
rect 179708 210294 179890 210354
rect 179708 210292 179714 210294
rect 19701 209674 19767 209677
rect 19701 209672 19810 209674
rect 19701 209616 19706 209672
rect 19762 209616 19810 209672
rect 19701 209611 19810 209616
rect 19750 209405 19810 209611
rect 19701 209400 19810 209405
rect 19701 209344 19706 209400
rect 19762 209344 19810 209400
rect 19701 209342 19810 209344
rect 19701 209339 19767 209342
rect 178401 205866 178467 205869
rect 178677 205866 178743 205869
rect 178401 205864 178743 205866
rect 178401 205808 178406 205864
rect 178462 205808 178682 205864
rect 178738 205808 178743 205864
rect 178401 205806 178743 205808
rect 178401 205803 178467 205806
rect 178677 205803 178743 205806
rect 179321 205866 179387 205869
rect 179454 205866 179460 205868
rect 179321 205864 179460 205866
rect 179321 205808 179326 205864
rect 179382 205808 179460 205864
rect 179321 205806 179460 205808
rect 179321 205803 179387 205806
rect 179454 205804 179460 205806
rect 179524 205804 179530 205868
rect 178166 205668 178172 205732
rect 178236 205730 178242 205732
rect 178236 205670 179706 205730
rect 178236 205668 178242 205670
rect 179646 205596 179706 205670
rect 179638 205532 179644 205596
rect 179708 205532 179714 205596
rect 583520 205580 584960 205820
rect 142061 203826 142127 203829
rect 143216 203826 143222 203828
rect 142061 203824 143222 203826
rect 142061 203768 142066 203824
rect 142122 203768 143222 203824
rect 142061 203766 143222 203768
rect 142061 203763 142127 203766
rect 143216 203764 143222 203766
rect 143286 203764 143292 203828
rect 179321 203826 179387 203829
rect 180006 203826 180012 203828
rect 179321 203824 180012 203826
rect 179321 203768 179326 203824
rect 179382 203768 180012 203824
rect 179321 203766 180012 203768
rect 179321 203763 179387 203766
rect 180006 203764 180012 203766
rect 180076 203764 180082 203828
rect 69749 203556 69815 203557
rect 71129 203556 71195 203557
rect 72233 203556 72299 203557
rect 73337 203556 73403 203557
rect 69749 203554 69782 203556
rect 69690 203552 69782 203554
rect 69690 203496 69754 203552
rect 69690 203494 69782 203496
rect 69749 203492 69782 203494
rect 69846 203492 69852 203556
rect 71129 203554 71142 203556
rect 71050 203552 71142 203554
rect 71050 203496 71134 203552
rect 71050 203494 71142 203496
rect 71129 203492 71142 203494
rect 71206 203492 71212 203556
rect 72224 203492 72230 203556
rect 72294 203554 72300 203556
rect 72294 203494 72386 203554
rect 72294 203492 72300 203494
rect 73312 203492 73318 203556
rect 73382 203554 73403 203556
rect 74349 203556 74415 203557
rect 75729 203556 75795 203557
rect 78029 203556 78095 203557
rect 229737 203556 229803 203557
rect 231117 203556 231183 203557
rect 232221 203556 232287 203557
rect 233325 203556 233391 203557
rect 234429 203556 234495 203557
rect 74349 203554 74406 203556
rect 73382 203552 73474 203554
rect 73398 203496 73474 203552
rect 73382 203494 73474 203496
rect 74314 203552 74406 203554
rect 74314 203496 74354 203552
rect 74314 203494 74406 203496
rect 73382 203492 73403 203494
rect 69749 203491 69815 203492
rect 71129 203491 71195 203492
rect 72233 203491 72299 203492
rect 73337 203491 73403 203492
rect 74349 203492 74406 203494
rect 74470 203492 74476 203556
rect 75729 203554 75766 203556
rect 75674 203552 75766 203554
rect 75674 203496 75734 203552
rect 75674 203494 75766 203496
rect 75729 203492 75766 203494
rect 75830 203492 75836 203556
rect 78029 203554 78078 203556
rect 77986 203552 78078 203554
rect 77986 203496 78034 203552
rect 77986 203494 78078 203496
rect 78029 203492 78078 203494
rect 78142 203492 78148 203556
rect 229737 203554 229782 203556
rect 229690 203552 229782 203554
rect 229690 203496 229742 203552
rect 229690 203494 229782 203496
rect 229737 203492 229782 203494
rect 229846 203492 229852 203556
rect 231117 203554 231142 203556
rect 231050 203552 231142 203554
rect 231050 203496 231122 203552
rect 231050 203494 231142 203496
rect 231117 203492 231142 203494
rect 231206 203492 231212 203556
rect 232221 203554 232230 203556
rect 232138 203552 232230 203554
rect 232138 203496 232226 203552
rect 232138 203494 232230 203496
rect 232221 203492 232230 203494
rect 232294 203492 232300 203556
rect 233312 203492 233318 203556
rect 233382 203554 233391 203556
rect 233382 203552 233474 203554
rect 233386 203496 233474 203552
rect 233382 203494 233474 203496
rect 233382 203492 233391 203494
rect 234400 203492 234406 203556
rect 234470 203554 234495 203556
rect 235717 203556 235783 203557
rect 237005 203556 237071 203557
rect 235717 203554 235766 203556
rect 234470 203552 234562 203554
rect 234490 203496 234562 203552
rect 234470 203494 234562 203496
rect 235674 203552 235766 203554
rect 235674 203496 235722 203552
rect 235674 203494 235766 203496
rect 234470 203492 234495 203494
rect 74349 203491 74415 203492
rect 75729 203491 75795 203492
rect 78029 203491 78095 203492
rect 229737 203491 229803 203492
rect 231117 203491 231183 203492
rect 232221 203491 232287 203492
rect 233325 203491 233391 203492
rect 234429 203491 234495 203492
rect 235717 203492 235766 203494
rect 235830 203492 235836 203556
rect 236984 203492 236990 203556
rect 237054 203554 237071 203556
rect 238017 203556 238083 203557
rect 238017 203554 238078 203556
rect 237054 203552 237146 203554
rect 237066 203496 237146 203552
rect 237054 203494 237146 203496
rect 237986 203552 238078 203554
rect 237986 203496 238022 203552
rect 237986 203494 238078 203496
rect 237054 203492 237071 203494
rect 235717 203491 235783 203492
rect 237005 203491 237071 203492
rect 238017 203492 238078 203494
rect 238142 203492 238148 203556
rect 238017 203491 238083 203492
rect 179638 203220 179644 203284
rect 179708 203282 179714 203284
rect 227478 203282 227484 203284
rect 179708 203222 227484 203282
rect 179708 203220 179714 203222
rect 227478 203220 227484 203222
rect 227548 203220 227554 203284
rect 178350 203084 178356 203148
rect 178420 203146 178426 203148
rect 226374 203146 226380 203148
rect 178420 203086 226380 203146
rect 178420 203084 178426 203086
rect 226374 203084 226380 203086
rect 226444 203084 226450 203148
rect 76925 203012 76991 203013
rect 76925 203010 76972 203012
rect 76880 203008 76972 203010
rect 76880 202952 76930 203008
rect 76880 202950 76972 202952
rect 76925 202948 76972 202950
rect 77036 202948 77042 203012
rect 179822 202948 179828 203012
rect 179892 203010 179898 203012
rect 228582 203010 228588 203012
rect 179892 202950 228588 203010
rect 179892 202948 179898 202950
rect 228582 202948 228588 202950
rect 228652 202948 228658 203012
rect 76925 202947 76991 202948
rect 19742 202812 19748 202876
rect 19812 202874 19818 202876
rect 47526 202874 47532 202876
rect 19812 202814 47532 202874
rect 19812 202812 19818 202814
rect 47526 202812 47532 202814
rect 47596 202812 47602 202876
rect 41597 202196 41663 202197
rect 41597 202194 41644 202196
rect 41552 202192 41644 202194
rect 41552 202136 41602 202192
rect 41552 202134 41644 202136
rect 41597 202132 41644 202134
rect 41708 202132 41714 202196
rect 41597 202131 41663 202132
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 35893 201380 35959 201381
rect 35893 201376 35940 201380
rect 36004 201378 36010 201380
rect 36537 201378 36603 201381
rect 37038 201378 37044 201380
rect 35893 201320 35898 201376
rect 35893 201316 35940 201320
rect 36004 201318 36050 201378
rect 36537 201376 37044 201378
rect 36537 201320 36542 201376
rect 36598 201320 37044 201376
rect 36537 201318 37044 201320
rect 36004 201316 36010 201318
rect 35893 201315 35959 201316
rect 36537 201315 36603 201318
rect 37038 201316 37044 201318
rect 37108 201316 37114 201380
rect 37273 201378 37339 201381
rect 38510 201378 38516 201380
rect 37273 201376 38516 201378
rect 37273 201320 37278 201376
rect 37334 201320 38516 201376
rect 37273 201318 38516 201320
rect 37273 201315 37339 201318
rect 38510 201316 38516 201318
rect 38580 201316 38586 201380
rect 38653 201378 38719 201381
rect 39614 201378 39620 201380
rect 38653 201376 39620 201378
rect 38653 201320 38658 201376
rect 38714 201320 39620 201376
rect 38653 201318 39620 201320
rect 38653 201315 38719 201318
rect 39614 201316 39620 201318
rect 39684 201316 39690 201380
rect 40033 201378 40099 201381
rect 44173 201380 44239 201381
rect 40534 201378 40540 201380
rect 40033 201376 40540 201378
rect 40033 201320 40038 201376
rect 40094 201320 40540 201376
rect 40033 201318 40540 201320
rect 40033 201315 40099 201318
rect 40534 201316 40540 201318
rect 40604 201316 40610 201380
rect 44173 201378 44220 201380
rect 44128 201376 44220 201378
rect 44128 201320 44178 201376
rect 44128 201318 44220 201320
rect 44173 201316 44220 201318
rect 44284 201316 44290 201380
rect 44357 201378 44423 201381
rect 44950 201378 44956 201380
rect 44357 201376 44956 201378
rect 44357 201320 44362 201376
rect 44418 201320 44956 201376
rect 44357 201318 44956 201320
rect 44173 201315 44239 201316
rect 44357 201315 44423 201318
rect 44950 201316 44956 201318
rect 45020 201316 45026 201380
rect 61694 201378 61700 201380
rect 45510 201318 61700 201378
rect 20662 201180 20668 201244
rect 20732 201242 20738 201244
rect 45510 201242 45570 201318
rect 61694 201316 61700 201318
rect 61764 201316 61770 201380
rect 63493 201378 63559 201381
rect 64086 201378 64092 201380
rect 63493 201376 64092 201378
rect 63493 201320 63498 201376
rect 63554 201320 64092 201376
rect 63493 201318 64092 201320
rect 63493 201315 63559 201318
rect 64086 201316 64092 201318
rect 64156 201316 64162 201380
rect 67633 201378 67699 201381
rect 68686 201378 68692 201380
rect 67633 201376 68692 201378
rect 67633 201320 67638 201376
rect 67694 201320 68692 201376
rect 67633 201318 68692 201320
rect 67633 201315 67699 201318
rect 68686 201316 68692 201318
rect 68756 201316 68762 201380
rect 79174 201316 79180 201380
rect 79244 201378 79250 201380
rect 79961 201378 80027 201381
rect 195973 201380 196039 201381
rect 195973 201378 196020 201380
rect 79244 201376 80027 201378
rect 79244 201320 79966 201376
rect 80022 201320 80027 201376
rect 79244 201318 80027 201320
rect 195928 201376 196020 201378
rect 195928 201320 195978 201376
rect 195928 201318 196020 201320
rect 79244 201316 79250 201318
rect 79961 201315 80027 201318
rect 195973 201316 196020 201318
rect 196084 201316 196090 201380
rect 196157 201378 196223 201381
rect 197118 201378 197124 201380
rect 196157 201376 197124 201378
rect 196157 201320 196162 201376
rect 196218 201320 197124 201376
rect 196157 201318 197124 201320
rect 195973 201315 196039 201316
rect 196157 201315 196223 201318
rect 197118 201316 197124 201318
rect 197188 201316 197194 201380
rect 197353 201378 197419 201381
rect 198222 201378 198228 201380
rect 197353 201376 198228 201378
rect 197353 201320 197358 201376
rect 197414 201320 198228 201376
rect 197353 201318 198228 201320
rect 197353 201315 197419 201318
rect 198222 201316 198228 201318
rect 198292 201316 198298 201380
rect 198733 201378 198799 201381
rect 199510 201378 199516 201380
rect 198733 201376 199516 201378
rect 198733 201320 198738 201376
rect 198794 201320 199516 201376
rect 198733 201318 199516 201320
rect 198733 201315 198799 201318
rect 199510 201316 199516 201318
rect 199580 201316 199586 201380
rect 200113 201378 200179 201381
rect 200614 201378 200620 201380
rect 200113 201376 200620 201378
rect 200113 201320 200118 201376
rect 200174 201320 200620 201376
rect 200113 201318 200620 201320
rect 200113 201315 200179 201318
rect 200614 201316 200620 201318
rect 200684 201316 200690 201380
rect 204345 201378 204411 201381
rect 205398 201378 205404 201380
rect 204345 201376 205404 201378
rect 204345 201320 204350 201376
rect 204406 201320 205404 201376
rect 204345 201318 205404 201320
rect 204345 201315 204411 201318
rect 205398 201316 205404 201318
rect 205468 201316 205474 201380
rect 211245 201378 211311 201381
rect 211654 201378 211660 201380
rect 211245 201376 211660 201378
rect 211245 201320 211250 201376
rect 211306 201320 211660 201376
rect 211245 201318 211660 201320
rect 211245 201315 211311 201318
rect 211654 201316 211660 201318
rect 211724 201316 211730 201380
rect 219985 201378 220051 201381
rect 220670 201378 220676 201380
rect 219985 201376 220676 201378
rect 219985 201320 219990 201376
rect 220046 201320 220676 201376
rect 219985 201318 220676 201320
rect 219985 201315 220051 201318
rect 220670 201316 220676 201318
rect 220740 201316 220746 201380
rect 222193 201378 222259 201381
rect 222878 201378 222884 201380
rect 222193 201376 222884 201378
rect 222193 201320 222198 201376
rect 222254 201320 222884 201376
rect 222193 201318 222884 201320
rect 222193 201315 222259 201318
rect 222878 201316 222884 201318
rect 222948 201316 222954 201380
rect 223573 201378 223639 201381
rect 224953 201380 225019 201381
rect 238937 201380 239003 201381
rect 303153 201380 303219 201381
rect 303521 201380 303587 201381
rect 223982 201378 223988 201380
rect 223573 201376 223988 201378
rect 223573 201320 223578 201376
rect 223634 201320 223988 201376
rect 223573 201318 223988 201320
rect 223573 201315 223639 201318
rect 223982 201316 223988 201318
rect 224052 201316 224058 201380
rect 224902 201316 224908 201380
rect 224972 201378 225019 201380
rect 238886 201378 238892 201380
rect 224972 201376 225064 201378
rect 225014 201320 225064 201376
rect 224972 201318 225064 201320
rect 238846 201318 238892 201378
rect 238956 201376 239003 201380
rect 303102 201378 303108 201380
rect 238998 201320 239003 201376
rect 224972 201316 225019 201318
rect 238886 201316 238892 201318
rect 238956 201316 239003 201320
rect 303062 201318 303108 201378
rect 303172 201376 303219 201380
rect 303214 201320 303219 201376
rect 303102 201316 303108 201318
rect 303172 201316 303219 201320
rect 303470 201316 303476 201380
rect 303540 201378 303587 201380
rect 303540 201376 303632 201378
rect 303582 201320 303632 201376
rect 303540 201318 303632 201320
rect 303540 201316 303587 201318
rect 224953 201315 225019 201316
rect 238937 201315 239003 201316
rect 303153 201315 303219 201316
rect 303521 201315 303587 201316
rect 20732 201182 45570 201242
rect 51073 201242 51139 201245
rect 51206 201242 51212 201244
rect 51073 201240 51212 201242
rect 51073 201184 51078 201240
rect 51134 201184 51212 201240
rect 51073 201182 51212 201184
rect 20732 201180 20738 201182
rect 51073 201179 51139 201182
rect 51206 201180 51212 201182
rect 51276 201180 51282 201244
rect 52453 201242 52519 201245
rect 55581 201244 55647 201245
rect 59353 201244 59419 201245
rect 53414 201242 53420 201244
rect 52453 201240 53420 201242
rect 52453 201184 52458 201240
rect 52514 201184 53420 201240
rect 52453 201182 53420 201184
rect 52453 201179 52519 201182
rect 53414 201180 53420 201182
rect 53484 201180 53490 201244
rect 55581 201242 55628 201244
rect 55536 201240 55628 201242
rect 55536 201184 55586 201240
rect 55536 201182 55628 201184
rect 55581 201180 55628 201182
rect 55692 201180 55698 201244
rect 59302 201180 59308 201244
rect 59372 201242 59419 201244
rect 62113 201242 62179 201245
rect 62798 201242 62804 201244
rect 59372 201240 59464 201242
rect 59414 201184 59464 201240
rect 59372 201182 59464 201184
rect 62113 201240 62804 201242
rect 62113 201184 62118 201240
rect 62174 201184 62804 201240
rect 62113 201182 62804 201184
rect 59372 201180 59419 201182
rect 55581 201179 55647 201180
rect 59353 201179 59419 201180
rect 62113 201179 62179 201182
rect 62798 201180 62804 201182
rect 62868 201180 62874 201244
rect 142061 201242 142127 201245
rect 143441 201242 143507 201245
rect 204253 201244 204319 201245
rect 142061 201240 143507 201242
rect 142061 201184 142066 201240
rect 142122 201184 143446 201240
rect 143502 201184 143507 201240
rect 142061 201182 143507 201184
rect 142061 201179 142127 201182
rect 143441 201179 143507 201182
rect 178534 201180 178540 201244
rect 178604 201242 178610 201244
rect 203006 201242 203012 201244
rect 178604 201182 203012 201242
rect 178604 201180 178610 201182
rect 203006 201180 203012 201182
rect 203076 201180 203082 201244
rect 204253 201242 204300 201244
rect 204208 201240 204300 201242
rect 204208 201184 204258 201240
rect 204208 201182 204300 201184
rect 204253 201180 204300 201182
rect 204364 201180 204370 201244
rect 214598 201242 214604 201244
rect 209730 201182 214604 201242
rect 204253 201179 204319 201180
rect 19006 201044 19012 201108
rect 19076 201106 19082 201108
rect 58014 201106 58020 201108
rect 19076 201046 58020 201106
rect 19076 201044 19082 201046
rect 58014 201044 58020 201046
rect 58084 201044 58090 201108
rect 59445 201106 59511 201109
rect 60590 201106 60596 201108
rect 59445 201104 60596 201106
rect 59445 201048 59450 201104
rect 59506 201048 60596 201104
rect 59445 201046 60596 201048
rect 59445 201043 59511 201046
rect 60590 201044 60596 201046
rect 60660 201044 60666 201108
rect 179454 201044 179460 201108
rect 179524 201106 179530 201108
rect 209730 201106 209790 201182
rect 214598 201180 214604 201182
rect 214668 201180 214674 201244
rect 215293 201242 215359 201245
rect 215886 201242 215892 201244
rect 215293 201240 215892 201242
rect 215293 201184 215298 201240
rect 215354 201184 215892 201240
rect 215293 201182 215892 201184
rect 215293 201179 215359 201182
rect 215886 201180 215892 201182
rect 215956 201180 215962 201244
rect 219433 201242 219499 201245
rect 219566 201242 219572 201244
rect 219433 201240 219572 201242
rect 219433 201184 219438 201240
rect 219494 201184 219572 201240
rect 219433 201182 219572 201184
rect 219433 201179 219499 201182
rect 219566 201180 219572 201182
rect 219636 201180 219642 201244
rect 179524 201046 209790 201106
rect 211153 201106 211219 201109
rect 212390 201106 212396 201108
rect 211153 201104 212396 201106
rect 211153 201048 211158 201104
rect 211214 201048 212396 201104
rect 211153 201046 212396 201048
rect 179524 201044 179530 201046
rect 211153 201043 211219 201046
rect 212390 201044 212396 201046
rect 212460 201044 212466 201108
rect 19190 200908 19196 200972
rect 19260 200970 19266 200972
rect 19260 200910 55230 200970
rect 19260 200908 19266 200910
rect 19558 200772 19564 200836
rect 19628 200834 19634 200836
rect 49693 200834 49759 200837
rect 50102 200834 50108 200836
rect 19628 200774 49618 200834
rect 19628 200772 19634 200774
rect 18638 200636 18644 200700
rect 18708 200698 18714 200700
rect 48630 200698 48636 200700
rect 18708 200638 48636 200698
rect 18708 200636 18714 200638
rect 48630 200636 48636 200638
rect 48700 200636 48706 200700
rect 49558 200698 49618 200774
rect 49693 200832 50108 200834
rect 49693 200776 49698 200832
rect 49754 200776 50108 200832
rect 49693 200774 50108 200776
rect 49693 200771 49759 200774
rect 50102 200772 50108 200774
rect 50172 200772 50178 200836
rect 51165 200834 51231 200837
rect 52310 200834 52316 200836
rect 51165 200832 52316 200834
rect 51165 200776 51170 200832
rect 51226 200776 52316 200832
rect 51165 200774 52316 200776
rect 51165 200771 51231 200774
rect 52310 200772 52316 200774
rect 52380 200772 52386 200836
rect 54518 200698 54524 200700
rect 49558 200638 54524 200698
rect 54518 200636 54524 200638
rect 54588 200636 54594 200700
rect 55170 200698 55230 200910
rect 180006 200908 180012 200972
rect 180076 200970 180082 200972
rect 213494 200970 213500 200972
rect 180076 200910 213500 200970
rect 180076 200908 180082 200910
rect 213494 200908 213500 200910
rect 213564 200908 213570 200972
rect 143441 200836 143507 200837
rect 143390 200772 143396 200836
rect 143460 200834 143507 200836
rect 143460 200832 143552 200834
rect 143502 200776 143552 200832
rect 143460 200774 143552 200776
rect 143460 200772 143507 200774
rect 179270 200772 179276 200836
rect 179340 200834 179346 200836
rect 208710 200834 208716 200836
rect 179340 200774 208716 200834
rect 179340 200772 179346 200774
rect 208710 200772 208716 200774
rect 208780 200772 208786 200836
rect 209865 200834 209931 200837
rect 209998 200834 210004 200836
rect 209865 200832 210004 200834
rect 209865 200776 209870 200832
rect 209926 200776 210004 200832
rect 209865 200774 210004 200776
rect 143441 200771 143507 200772
rect 209865 200771 209931 200774
rect 209998 200772 210004 200774
rect 210068 200772 210074 200836
rect 56910 200698 56916 200700
rect 55170 200638 56916 200698
rect 56910 200636 56916 200638
rect 56980 200636 56986 200700
rect 62021 200698 62087 200701
rect 352557 200698 352623 200701
rect 62021 200696 352623 200698
rect 62021 200640 62026 200696
rect 62082 200640 352562 200696
rect 352618 200640 352623 200696
rect 62021 200638 352623 200640
rect 62021 200635 62087 200638
rect 352557 200635 352623 200638
rect 19374 200500 19380 200564
rect 19444 200562 19450 200564
rect 67766 200562 67772 200564
rect 19444 200502 67772 200562
rect 19444 200500 19450 200502
rect 67766 200500 67772 200502
rect 67836 200500 67842 200564
rect 178902 200500 178908 200564
rect 178972 200562 178978 200564
rect 201309 200562 201375 200565
rect 178972 200560 201375 200562
rect 178972 200504 201314 200560
rect 201370 200504 201375 200560
rect 178972 200502 201375 200504
rect 178972 200500 178978 200502
rect 201309 200499 201375 200502
rect 201493 200562 201559 200565
rect 201718 200562 201724 200564
rect 201493 200560 201724 200562
rect 201493 200504 201498 200560
rect 201554 200504 201724 200560
rect 201493 200502 201724 200504
rect 201493 200499 201559 200502
rect 201718 200500 201724 200502
rect 201788 200500 201794 200564
rect 201861 200562 201927 200565
rect 207054 200562 207060 200564
rect 201861 200560 207060 200562
rect 201861 200504 201866 200560
rect 201922 200504 207060 200560
rect 201861 200502 207060 200504
rect 201861 200499 201927 200502
rect 207054 200500 207060 200502
rect 207124 200500 207130 200564
rect 66253 200428 66319 200429
rect 18822 200364 18828 200428
rect 18892 200426 18898 200428
rect 43110 200426 43116 200428
rect 18892 200366 43116 200426
rect 18892 200364 18898 200366
rect 43110 200364 43116 200366
rect 43180 200364 43186 200428
rect 66253 200426 66300 200428
rect 66208 200424 66300 200426
rect 66208 200368 66258 200424
rect 66208 200366 66300 200368
rect 66253 200364 66300 200366
rect 66364 200364 66370 200428
rect 178953 200426 179019 200429
rect 218646 200426 218652 200428
rect 178953 200424 218652 200426
rect 178953 200368 178958 200424
rect 179014 200368 218652 200424
rect 178953 200366 218652 200368
rect 66253 200363 66319 200364
rect 178953 200363 179019 200366
rect 218646 200364 218652 200366
rect 218716 200364 218722 200428
rect 18454 200228 18460 200292
rect 18524 200290 18530 200292
rect 46422 200290 46428 200292
rect 18524 200230 46428 200290
rect 18524 200228 18530 200230
rect 46422 200228 46428 200230
rect 46492 200228 46498 200292
rect 64638 200228 64644 200292
rect 64708 200290 64714 200292
rect 64873 200290 64939 200293
rect 64708 200288 64939 200290
rect 64708 200232 64878 200288
rect 64934 200232 64939 200288
rect 64708 200230 64939 200232
rect 64708 200228 64714 200230
rect 64873 200227 64939 200230
rect 178718 200228 178724 200292
rect 178788 200290 178794 200292
rect 216990 200290 216996 200292
rect 178788 200230 216996 200290
rect 178788 200228 178794 200230
rect 216990 200228 216996 200230
rect 217060 200228 217066 200292
rect 220813 200290 220879 200293
rect 221222 200290 221228 200292
rect 220813 200288 221228 200290
rect 220813 200232 220818 200288
rect 220874 200232 221228 200288
rect 220813 200230 221228 200232
rect 220813 200227 220879 200230
rect 221222 200228 221228 200230
rect 221292 200228 221298 200292
rect 179086 200092 179092 200156
rect 179156 200154 179162 200156
rect 201125 200154 201191 200157
rect 179156 200152 201191 200154
rect 179156 200096 201130 200152
rect 201186 200096 201191 200152
rect 179156 200094 201191 200096
rect 179156 200092 179162 200094
rect 201125 200091 201191 200094
rect 201309 200154 201375 200157
rect 206502 200154 206508 200156
rect 201309 200152 206508 200154
rect 201309 200096 201314 200152
rect 201370 200096 206508 200152
rect 201309 200094 206508 200096
rect 201309 200091 201375 200094
rect 206502 200092 206508 200094
rect 206572 200092 206578 200156
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 213500 408444 213564 408508
rect 216260 408444 216324 408508
rect 226196 408504 226260 408508
rect 226196 408448 226246 408504
rect 226246 408448 226260 408504
rect 226196 408444 226260 408448
rect 228588 408444 228652 408508
rect 251036 408504 251100 408508
rect 251036 408448 251086 408504
rect 251086 408448 251100 408504
rect 251036 408444 251100 408448
rect 253612 408444 253676 408508
rect 258580 408444 258644 408508
rect 263548 408444 263612 408508
rect 265940 408444 266004 408508
rect 273668 408444 273732 408508
rect 278452 408444 278516 408508
rect 221044 408308 221108 408372
rect 223436 408368 223500 408372
rect 223436 408312 223486 408368
rect 223486 408312 223500 408368
rect 223436 408308 223500 408312
rect 271092 408308 271156 408372
rect 286180 408308 286244 408372
rect 90956 408172 91020 408236
rect 268516 408036 268580 408100
rect 139716 407900 139780 407964
rect 71084 407764 71148 407828
rect 93532 407764 93596 407828
rect 66116 407688 66180 407692
rect 66116 407632 66166 407688
rect 66166 407632 66180 407688
rect 66116 407628 66180 407632
rect 101076 407628 101140 407692
rect 106044 407492 106108 407556
rect 103652 407356 103716 407420
rect 63540 407220 63604 407284
rect 68508 407220 68572 407284
rect 51028 407084 51092 407148
rect 56180 407084 56244 407148
rect 58572 407084 58636 407148
rect 98684 407084 98748 407148
rect 108436 407084 108500 407148
rect 111012 407084 111076 407148
rect 113588 407084 113652 407148
rect 115980 407084 116044 407148
rect 118556 407144 118620 407148
rect 118556 407088 118606 407144
rect 118606 407088 118620 407144
rect 118556 407084 118620 407088
rect 121132 407084 121196 407148
rect 123340 407084 123404 407148
rect 126100 407084 126164 407148
rect 138428 407084 138492 407148
rect 150940 407084 151004 407148
rect 208716 407084 208780 407148
rect 211108 407144 211172 407148
rect 211108 407088 211122 407144
rect 211122 407088 211172 407144
rect 211108 407084 211172 407088
rect 218468 407084 218532 407148
rect 231164 407084 231228 407148
rect 233556 407084 233620 407148
rect 236132 407084 236196 407148
rect 240916 407084 240980 407148
rect 246068 407084 246132 407148
rect 248644 407084 248708 407148
rect 256004 407084 256068 407148
rect 261156 407084 261220 407148
rect 276060 407084 276124 407148
rect 283420 407084 283484 407148
rect 298508 407084 298572 407148
rect 299796 407084 299860 407148
rect 310836 407084 310900 407148
rect 78444 406540 78508 406604
rect 81020 406464 81084 406468
rect 81020 406408 81070 406464
rect 81070 406408 81084 406464
rect 81020 406404 81084 406408
rect 83596 406464 83660 406468
rect 86172 406600 86236 406604
rect 86172 406544 86222 406600
rect 86222 406544 86236 406600
rect 86172 406540 86236 406544
rect 88564 406600 88628 406604
rect 88564 406544 88614 406600
rect 88614 406544 88628 406600
rect 88564 406540 88628 406544
rect 95924 406600 95988 406604
rect 95924 406544 95974 406600
rect 95974 406544 95988 406600
rect 95924 406540 95988 406544
rect 238524 406600 238588 406604
rect 238524 406544 238574 406600
rect 238574 406544 238588 406600
rect 238524 406540 238588 406544
rect 243676 406600 243740 406604
rect 243676 406544 243726 406600
rect 243726 406544 243740 406600
rect 243676 406540 243740 406544
rect 281028 406600 281092 406604
rect 281028 406544 281078 406600
rect 281078 406544 281092 406600
rect 281028 406540 281092 406544
rect 83596 406408 83646 406464
rect 83646 406408 83660 406464
rect 83596 406404 83660 406408
rect 48702 406192 48766 406196
rect 48702 406136 48742 406192
rect 48742 406136 48766 406192
rect 48702 406132 48766 406136
rect 53462 406192 53526 406196
rect 53462 406136 53470 406192
rect 53470 406136 53526 406192
rect 53462 406132 53526 406136
rect 61078 406192 61142 406196
rect 61078 406136 61106 406192
rect 61106 406136 61142 406192
rect 61078 406132 61142 406136
rect 73590 406132 73654 406196
rect 76174 406132 76238 406196
rect 143358 322008 143422 322012
rect 143358 321952 143410 322008
rect 143410 321952 143422 322008
rect 143358 321948 143422 321952
rect 226932 321948 226996 322012
rect 227606 321948 227670 322012
rect 228694 321948 228758 322012
rect 68692 321812 68756 321876
rect 179644 321812 179708 321876
rect 66484 321676 66548 321740
rect 179460 321736 179524 321740
rect 179460 321680 179474 321736
rect 179474 321680 179524 321736
rect 179460 321676 179524 321680
rect 226380 321736 226444 321740
rect 226380 321680 226394 321736
rect 226394 321680 226444 321736
rect 226380 321676 226444 321680
rect 62804 321600 62868 321604
rect 62804 321544 62818 321600
rect 62818 321544 62868 321600
rect 62804 321540 62868 321544
rect 63908 321600 63972 321604
rect 63908 321544 63922 321600
rect 63922 321544 63972 321600
rect 63908 321540 63972 321544
rect 67588 321600 67652 321604
rect 67588 321544 67638 321600
rect 67638 321544 67652 321600
rect 67588 321540 67652 321544
rect 180012 321540 180076 321604
rect 19012 321404 19076 321468
rect 58204 321404 58268 321468
rect 219204 321404 219268 321468
rect 220676 321404 220740 321468
rect 19196 321268 19260 321332
rect 56916 321268 56980 321332
rect 54524 321132 54588 321196
rect 19380 320588 19444 320652
rect 61700 320588 61764 320652
rect 207612 320588 207676 320652
rect 221780 320648 221844 320652
rect 221780 320592 221830 320648
rect 221830 320592 221844 320648
rect 221780 320588 221844 320592
rect 20668 320452 20732 320516
rect 74580 320512 74644 320516
rect 74580 320456 74630 320512
rect 74630 320456 74644 320512
rect 74580 320452 74644 320456
rect 143212 320512 143276 320516
rect 143212 320456 143262 320512
rect 143262 320456 143276 320512
rect 143212 320452 143276 320456
rect 43116 320180 43180 320244
rect 178540 320240 178604 320244
rect 178540 320184 178590 320240
rect 178590 320184 178604 320240
rect 178540 320180 178604 320184
rect 178724 320240 178788 320244
rect 178724 320184 178774 320240
rect 178774 320184 178788 320240
rect 178724 320180 178788 320184
rect 179828 320180 179892 320244
rect 44220 320104 44284 320108
rect 44220 320048 44234 320104
rect 44234 320048 44284 320104
rect 18828 319772 18892 319836
rect 44220 320044 44284 320048
rect 44956 320104 45020 320108
rect 44956 320048 45006 320104
rect 45006 320048 45020 320104
rect 44956 320044 45020 320048
rect 50108 320104 50172 320108
rect 50108 320048 50158 320104
rect 50158 320048 50172 320104
rect 50108 320044 50172 320048
rect 51212 320104 51276 320108
rect 51212 320048 51262 320104
rect 51262 320048 51276 320104
rect 51212 320044 51276 320048
rect 52316 320104 52380 320108
rect 52316 320048 52366 320104
rect 52366 320048 52380 320104
rect 52316 320044 52380 320048
rect 53420 320104 53484 320108
rect 53420 320048 53470 320104
rect 53470 320048 53484 320104
rect 53420 320044 53484 320048
rect 59308 320104 59372 320108
rect 59308 320048 59358 320104
rect 59358 320048 59372 320104
rect 59308 320044 59372 320048
rect 65380 320104 65444 320108
rect 65380 320048 65394 320104
rect 65394 320048 65444 320104
rect 65380 320044 65444 320048
rect 68692 320104 68756 320108
rect 68692 320048 68706 320104
rect 68706 320048 68756 320104
rect 68692 320044 68756 320048
rect 71084 320104 71148 320108
rect 71084 320048 71134 320104
rect 71134 320048 71148 320104
rect 71084 320044 71148 320048
rect 72188 320104 72252 320108
rect 72188 320048 72202 320104
rect 72202 320048 72252 320104
rect 72188 320044 72252 320048
rect 73292 320104 73356 320108
rect 73292 320048 73342 320104
rect 73342 320048 73356 320104
rect 73292 320044 73356 320048
rect 75684 320104 75748 320108
rect 75684 320048 75734 320104
rect 75734 320048 75748 320104
rect 75684 320044 75748 320048
rect 79180 320104 79244 320108
rect 79180 320048 79230 320104
rect 79230 320048 79244 320104
rect 79180 320044 79244 320048
rect 200620 320044 200684 320108
rect 203196 320104 203260 320108
rect 203196 320048 203210 320104
rect 203210 320048 203260 320104
rect 203196 320044 203260 320048
rect 204300 320104 204364 320108
rect 204300 320048 204350 320104
rect 204350 320048 204364 320104
rect 204300 320044 204364 320048
rect 211660 320044 211724 320108
rect 223988 320044 224052 320108
rect 226380 320044 226444 320108
rect 231164 320104 231228 320108
rect 231164 320048 231214 320104
rect 231214 320048 231228 320104
rect 231164 320044 231228 320048
rect 36124 319968 36188 319972
rect 36124 319912 36138 319968
rect 36138 319912 36188 319968
rect 36124 319908 36188 319912
rect 39620 319968 39684 319972
rect 39620 319912 39634 319968
rect 39634 319912 39684 319968
rect 39620 319908 39684 319912
rect 60596 319908 60660 319972
rect 66484 319968 66548 319972
rect 66484 319912 66498 319968
rect 66498 319912 66548 319968
rect 66484 319908 66548 319912
rect 214604 319908 214668 319972
rect 226932 319968 226996 319972
rect 226932 319912 226982 319968
rect 226982 319912 226996 319968
rect 226932 319908 226996 319912
rect 229692 319908 229756 319972
rect 210004 319772 210068 319836
rect 55628 319636 55692 319700
rect 78260 319636 78324 319700
rect 215892 319636 215956 319700
rect 216996 319636 217060 319700
rect 218652 319636 218716 319700
rect 232268 319636 232332 319700
rect 18644 319500 18708 319564
rect 48636 319500 48700 319564
rect 179276 319500 179340 319564
rect 19564 319364 19628 319428
rect 47532 319364 47596 319428
rect 179092 319364 179156 319428
rect 40540 319228 40604 319292
rect 42380 319228 42444 319292
rect 69796 319228 69860 319292
rect 76972 319228 77036 319292
rect 236868 319500 236932 319564
rect 196020 319424 196084 319428
rect 196020 319368 196070 319424
rect 196070 319368 196084 319424
rect 196020 319364 196084 319368
rect 198228 319364 198292 319428
rect 199516 319364 199580 319428
rect 201724 319228 201788 319292
rect 213500 319364 213564 319428
rect 222884 319424 222948 319428
rect 222884 319368 222898 319424
rect 222898 319368 222948 319424
rect 222884 319364 222948 319368
rect 303108 319424 303172 319428
rect 303108 319368 303122 319424
rect 303122 319368 303172 319424
rect 303108 319364 303172 319368
rect 37044 319092 37108 319156
rect 38516 319092 38580 319156
rect 46428 319092 46492 319156
rect 177988 319092 178052 319156
rect 178908 319092 178972 319156
rect 206508 319228 206572 319292
rect 208716 319228 208780 319292
rect 224908 319228 224972 319292
rect 234292 319228 234356 319292
rect 235580 319228 235644 319292
rect 303476 319228 303540 319292
rect 205404 319092 205468 319156
rect 212396 319092 212460 319156
rect 237972 319152 238036 319156
rect 237972 319096 238022 319152
rect 238022 319096 238036 319152
rect 237972 319092 238036 319096
rect 239076 318956 239140 319020
rect 177988 318820 178052 318884
rect 180564 318880 180628 318884
rect 180564 318824 180578 318880
rect 180578 318824 180628 318880
rect 180564 318820 180628 318824
rect 197124 318820 197188 318884
rect 233372 318820 233436 318884
rect 19564 316236 19628 316300
rect 19564 316100 19628 316164
rect 19380 315964 19444 316028
rect 19380 315828 19444 315892
rect 20668 315828 20732 315892
rect 19380 306580 19444 306644
rect 19380 306444 19444 306508
rect 20852 306444 20916 306508
rect 19380 306308 19444 306372
rect 20852 306308 20916 306372
rect 19380 306172 19444 306236
rect 19380 296924 19444 296988
rect 19380 296788 19444 296852
rect 20668 296788 20732 296852
rect 19380 296652 19444 296716
rect 19380 296516 19444 296580
rect 20668 296516 20732 296580
rect 48636 291076 48700 291140
rect 51028 291076 51092 291140
rect 53420 291076 53484 291140
rect 56548 291136 56612 291140
rect 56548 291080 56562 291136
rect 56562 291080 56612 291136
rect 56548 291076 56612 291080
rect 58572 291076 58636 291140
rect 61148 291076 61212 291140
rect 64092 291076 64156 291140
rect 68508 291076 68572 291140
rect 71084 291076 71148 291140
rect 76236 291076 76300 291140
rect 78444 291076 78508 291140
rect 81020 291076 81084 291140
rect 83596 291076 83660 291140
rect 86172 291076 86236 291140
rect 88564 291076 88628 291140
rect 90956 291136 91020 291140
rect 90956 291080 91006 291136
rect 91006 291080 91020 291136
rect 90956 291076 91020 291080
rect 93532 291076 93596 291140
rect 98684 291076 98748 291140
rect 106044 291076 106108 291140
rect 115980 291076 116044 291140
rect 208716 291076 208780 291140
rect 210740 291076 210804 291140
rect 213500 291076 213564 291140
rect 216260 291076 216324 291140
rect 218652 291076 218716 291140
rect 221044 291076 221108 291140
rect 223436 291136 223500 291140
rect 223436 291080 223486 291136
rect 223486 291080 223500 291136
rect 223436 291076 223500 291080
rect 226196 291136 226260 291140
rect 226196 291080 226246 291136
rect 226246 291080 226260 291136
rect 226196 291076 226260 291080
rect 228588 291076 228652 291140
rect 231164 291076 231228 291140
rect 238524 291076 238588 291140
rect 240916 291076 240980 291140
rect 244044 291076 244108 291140
rect 246068 291076 246132 291140
rect 248644 291076 248708 291140
rect 251036 291136 251100 291140
rect 251036 291080 251086 291136
rect 251086 291080 251100 291136
rect 251036 291076 251100 291080
rect 253612 291076 253676 291140
rect 256004 291076 256068 291140
rect 258580 291076 258644 291140
rect 263548 291076 263612 291140
rect 268516 291076 268580 291140
rect 271092 291076 271156 291140
rect 273668 291076 273732 291140
rect 276244 291076 276308 291140
rect 281028 291076 281092 291140
rect 283788 291076 283852 291140
rect 101076 290940 101140 291004
rect 113220 290940 113284 291004
rect 236500 290940 236564 291004
rect 111012 290804 111076 290868
rect 139716 290804 139780 290868
rect 64828 290668 64892 290732
rect 103836 290668 103900 290732
rect 118556 290728 118620 290732
rect 118556 290672 118606 290728
rect 118606 290672 118620 290728
rect 118556 290668 118620 290672
rect 265940 290668 266004 290732
rect 277348 290668 277412 290732
rect 126100 290396 126164 290460
rect 138428 290396 138492 290460
rect 260972 290396 261036 290460
rect 73476 290260 73540 290324
rect 120764 290260 120828 290324
rect 96292 290124 96356 290188
rect 108436 289988 108500 290052
rect 122788 290048 122852 290052
rect 122788 289992 122838 290048
rect 122838 289992 122852 290048
rect 122788 289988 122852 289992
rect 233556 289988 233620 290052
rect 286180 289852 286244 289916
rect 298508 289852 298572 289916
rect 299612 289912 299676 289916
rect 299612 289856 299662 289912
rect 299662 289856 299676 289912
rect 299612 289852 299676 289856
rect 310836 289912 310900 289916
rect 310836 289856 310850 289912
rect 310850 289856 310900 289912
rect 310836 289852 310900 289856
rect 19380 288900 19444 288964
rect 19748 288900 19812 288964
rect 178356 288764 178420 288828
rect 179276 288764 179340 288828
rect 19380 288492 19444 288556
rect 20852 288492 20916 288556
rect 179276 287812 179340 287876
rect 179644 287812 179708 287876
rect 18460 287676 18524 287740
rect 179644 287676 179708 287740
rect 180012 287676 180076 287740
rect 150838 287464 150902 287468
rect 150838 287408 150898 287464
rect 150898 287408 150902 287464
rect 150838 287404 150902 287408
rect 180564 287404 180628 287468
rect 178172 267684 178236 267748
rect 178172 258164 178236 258228
rect 178172 257892 178236 257956
rect 178172 253812 178236 253876
rect 179828 245924 179892 245988
rect 179828 245652 179892 245716
rect 179644 244700 179708 244764
rect 179276 244564 179340 244628
rect 178356 244292 178420 244356
rect 179276 244292 179340 244356
rect 179644 244292 179708 244356
rect 179644 243944 179708 243948
rect 179644 243888 179658 243944
rect 179658 243888 179708 243944
rect 179644 243884 179708 243888
rect 179828 243884 179892 243948
rect 179644 243748 179708 243812
rect 179828 243612 179892 243676
rect 178356 239396 178420 239460
rect 179276 239396 179340 239460
rect 179276 236540 179340 236604
rect 179644 236540 179708 236604
rect 179644 236464 179708 236468
rect 179644 236408 179658 236464
rect 179658 236408 179708 236464
rect 179644 236404 179708 236408
rect 179276 234772 179340 234836
rect 179276 234636 179340 234700
rect 178172 234364 178236 234428
rect 179276 234364 179340 234428
rect 179276 234228 179340 234292
rect 179460 233004 179524 233068
rect 179644 233004 179708 233068
rect 179828 233004 179892 233068
rect 179460 232732 179524 232796
rect 179644 232732 179708 232796
rect 179828 232732 179892 232796
rect 178172 224844 178236 224908
rect 179460 224844 179524 224908
rect 179644 224844 179708 224908
rect 177988 224708 178052 224772
rect 179460 224708 179524 224772
rect 179644 224572 179708 224636
rect 177804 222668 177868 222732
rect 179276 222668 179340 222732
rect 178356 220084 178420 220148
rect 179276 220084 179340 220148
rect 179828 210564 179892 210628
rect 179644 210292 179708 210356
rect 179460 205804 179524 205868
rect 178172 205668 178236 205732
rect 179644 205532 179708 205596
rect 143222 203764 143286 203828
rect 180012 203764 180076 203828
rect 69782 203552 69846 203556
rect 69782 203496 69810 203552
rect 69810 203496 69846 203552
rect 69782 203492 69846 203496
rect 71142 203552 71206 203556
rect 71142 203496 71190 203552
rect 71190 203496 71206 203552
rect 71142 203492 71206 203496
rect 72230 203552 72294 203556
rect 72230 203496 72238 203552
rect 72238 203496 72294 203552
rect 72230 203492 72294 203496
rect 73318 203552 73382 203556
rect 73318 203496 73342 203552
rect 73342 203496 73382 203552
rect 73318 203492 73382 203496
rect 74406 203552 74470 203556
rect 74406 203496 74410 203552
rect 74410 203496 74470 203552
rect 74406 203492 74470 203496
rect 75766 203552 75830 203556
rect 75766 203496 75790 203552
rect 75790 203496 75830 203552
rect 75766 203492 75830 203496
rect 78078 203552 78142 203556
rect 78078 203496 78090 203552
rect 78090 203496 78142 203552
rect 78078 203492 78142 203496
rect 229782 203552 229846 203556
rect 229782 203496 229798 203552
rect 229798 203496 229846 203552
rect 229782 203492 229846 203496
rect 231142 203552 231206 203556
rect 231142 203496 231178 203552
rect 231178 203496 231206 203552
rect 231142 203492 231206 203496
rect 232230 203552 232294 203556
rect 232230 203496 232282 203552
rect 232282 203496 232294 203552
rect 232230 203492 232294 203496
rect 233318 203552 233382 203556
rect 233318 203496 233330 203552
rect 233330 203496 233382 203552
rect 233318 203492 233382 203496
rect 234406 203552 234470 203556
rect 234406 203496 234434 203552
rect 234434 203496 234470 203552
rect 234406 203492 234470 203496
rect 235766 203552 235830 203556
rect 235766 203496 235778 203552
rect 235778 203496 235830 203552
rect 235766 203492 235830 203496
rect 236990 203552 237054 203556
rect 236990 203496 237010 203552
rect 237010 203496 237054 203552
rect 236990 203492 237054 203496
rect 238078 203492 238142 203556
rect 179644 203220 179708 203284
rect 227484 203220 227548 203284
rect 178356 203084 178420 203148
rect 226380 203084 226444 203148
rect 76972 203008 77036 203012
rect 76972 202952 76986 203008
rect 76986 202952 77036 203008
rect 76972 202948 77036 202952
rect 179828 202948 179892 203012
rect 228588 202948 228652 203012
rect 19748 202812 19812 202876
rect 47532 202812 47596 202876
rect 41644 202192 41708 202196
rect 41644 202136 41658 202192
rect 41658 202136 41708 202192
rect 41644 202132 41708 202136
rect 35940 201376 36004 201380
rect 35940 201320 35954 201376
rect 35954 201320 36004 201376
rect 35940 201316 36004 201320
rect 37044 201316 37108 201380
rect 38516 201316 38580 201380
rect 39620 201316 39684 201380
rect 40540 201316 40604 201380
rect 44220 201376 44284 201380
rect 44220 201320 44234 201376
rect 44234 201320 44284 201376
rect 44220 201316 44284 201320
rect 44956 201316 45020 201380
rect 20668 201180 20732 201244
rect 61700 201316 61764 201380
rect 64092 201316 64156 201380
rect 68692 201316 68756 201380
rect 79180 201316 79244 201380
rect 196020 201376 196084 201380
rect 196020 201320 196034 201376
rect 196034 201320 196084 201376
rect 196020 201316 196084 201320
rect 197124 201316 197188 201380
rect 198228 201316 198292 201380
rect 199516 201316 199580 201380
rect 200620 201316 200684 201380
rect 205404 201316 205468 201380
rect 211660 201316 211724 201380
rect 220676 201316 220740 201380
rect 222884 201316 222948 201380
rect 223988 201316 224052 201380
rect 224908 201376 224972 201380
rect 224908 201320 224958 201376
rect 224958 201320 224972 201376
rect 224908 201316 224972 201320
rect 238892 201376 238956 201380
rect 238892 201320 238942 201376
rect 238942 201320 238956 201376
rect 238892 201316 238956 201320
rect 303108 201376 303172 201380
rect 303108 201320 303158 201376
rect 303158 201320 303172 201376
rect 303108 201316 303172 201320
rect 303476 201376 303540 201380
rect 303476 201320 303526 201376
rect 303526 201320 303540 201376
rect 303476 201316 303540 201320
rect 51212 201180 51276 201244
rect 53420 201180 53484 201244
rect 55628 201240 55692 201244
rect 55628 201184 55642 201240
rect 55642 201184 55692 201240
rect 55628 201180 55692 201184
rect 59308 201240 59372 201244
rect 59308 201184 59358 201240
rect 59358 201184 59372 201240
rect 59308 201180 59372 201184
rect 62804 201180 62868 201244
rect 178540 201180 178604 201244
rect 203012 201180 203076 201244
rect 204300 201240 204364 201244
rect 204300 201184 204314 201240
rect 204314 201184 204364 201240
rect 204300 201180 204364 201184
rect 19012 201044 19076 201108
rect 58020 201044 58084 201108
rect 60596 201044 60660 201108
rect 179460 201044 179524 201108
rect 214604 201180 214668 201244
rect 215892 201180 215956 201244
rect 219572 201180 219636 201244
rect 212396 201044 212460 201108
rect 19196 200908 19260 200972
rect 19564 200772 19628 200836
rect 18644 200636 18708 200700
rect 48636 200636 48700 200700
rect 50108 200772 50172 200836
rect 52316 200772 52380 200836
rect 54524 200636 54588 200700
rect 180012 200908 180076 200972
rect 213500 200908 213564 200972
rect 143396 200832 143460 200836
rect 143396 200776 143446 200832
rect 143446 200776 143460 200832
rect 143396 200772 143460 200776
rect 179276 200772 179340 200836
rect 208716 200772 208780 200836
rect 210004 200772 210068 200836
rect 56916 200636 56980 200700
rect 19380 200500 19444 200564
rect 67772 200500 67836 200564
rect 178908 200500 178972 200564
rect 201724 200500 201788 200564
rect 207060 200500 207124 200564
rect 18828 200364 18892 200428
rect 43116 200364 43180 200428
rect 66300 200424 66364 200428
rect 66300 200368 66314 200424
rect 66314 200368 66364 200424
rect 66300 200364 66364 200368
rect 218652 200364 218716 200428
rect 18460 200228 18524 200292
rect 46428 200228 46492 200292
rect 64644 200228 64708 200292
rect 178724 200228 178788 200292
rect 216996 200228 217060 200292
rect 221228 200228 221292 200292
rect 179092 200092 179156 200156
rect 206508 200092 206572 200156
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 3739 371380 3805 371381
rect 3739 371316 3740 371380
rect 3804 371316 3805 371380
rect 3739 371315 3805 371316
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 3555 358460 3621 358461
rect 3555 358396 3556 358460
rect 3620 358396 3621 358460
rect 3555 358395 3621 358396
rect 3371 345404 3437 345405
rect 3371 345340 3372 345404
rect 3436 345340 3437 345404
rect 3371 345339 3437 345340
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 3374 315893 3434 345339
rect 3558 330309 3618 358395
rect 3742 344725 3802 371315
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 3739 344724 3805 344725
rect 3739 344660 3740 344724
rect 3804 344660 3805 344724
rect 3739 344659 3805 344660
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 3555 330308 3621 330309
rect 3555 330244 3556 330308
rect 3620 330244 3621 330308
rect 3555 330243 3621 330244
rect 3739 319292 3805 319293
rect 3739 319228 3740 319292
rect 3804 319228 3805 319292
rect 3739 319227 3805 319228
rect 3371 315892 3437 315893
rect 3371 315828 3372 315892
rect 3436 315828 3437 315892
rect 3371 315827 3437 315828
rect 3555 306236 3621 306237
rect 3555 306172 3556 306236
rect 3620 306172 3621 306236
rect 3555 306171 3621 306172
rect 3371 293180 3437 293181
rect 3371 293116 3372 293180
rect 3436 293116 3437 293180
rect 3371 293115 3437 293116
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 3374 272645 3434 293115
rect 3558 287061 3618 306171
rect 3742 301477 3802 319227
rect 3739 301476 3805 301477
rect 3739 301412 3740 301476
rect 3804 301412 3805 301476
rect 3739 301411 3805 301412
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 3555 287060 3621 287061
rect 3555 286996 3556 287060
rect 3620 286996 3621 287060
rect 3555 286995 3621 286996
rect 3371 272644 3437 272645
rect 3371 272580 3372 272644
rect 3436 272580 3437 272644
rect 3371 272579 3437 272580
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 5514 259174 6134 294618
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 8155 267204 8221 267205
rect 8155 267140 8156 267204
rect 8220 267140 8221 267204
rect 8155 267139 8221 267140
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 8158 258229 8218 267139
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 8155 258228 8221 258229
rect 8155 258164 8156 258228
rect 8220 258164 8221 258228
rect 8155 258163 8221 258164
rect 7419 254148 7485 254149
rect 7419 254084 7420 254148
rect 7484 254084 7485 254148
rect 7419 254083 7485 254084
rect 7422 243813 7482 254083
rect 7419 243812 7485 243813
rect 7419 243748 7420 243812
rect 7484 243748 7485 243812
rect 7419 243747 7485 243748
rect 7419 241092 7485 241093
rect 7419 241028 7420 241092
rect 7484 241028 7485 241092
rect 7419 241027 7485 241028
rect 7422 229397 7482 241027
rect 7419 229396 7485 229397
rect 7419 229332 7420 229396
rect 7484 229332 7485 229396
rect 7419 229331 7485 229332
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 6315 188868 6381 188869
rect 6315 188804 6316 188868
rect 6380 188804 6381 188868
rect 6315 188803 6381 188804
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 6318 186149 6378 188803
rect 6315 186148 6381 186149
rect 6315 186084 6316 186148
rect 6380 186084 6381 186148
rect 6315 186083 6381 186084
rect 6315 171732 6381 171733
rect 6315 171668 6316 171732
rect 6380 171668 6381 171732
rect 6315 171667 6381 171668
rect 6318 162893 6378 171667
rect 6315 162892 6381 162893
rect 6315 162828 6316 162892
rect 6380 162828 6381 162892
rect 6315 162827 6381 162828
rect 6315 157316 6381 157317
rect 6315 157252 6316 157316
rect 6380 157252 6381 157316
rect 6315 157251 6381 157252
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 4843 142900 4909 142901
rect 4843 142836 4844 142900
rect 4908 142836 4909 142900
rect 4843 142835 4909 142836
rect 4846 136781 4906 142835
rect 4843 136780 4909 136781
rect 4843 136716 4844 136780
rect 4908 136716 4909 136780
rect 4843 136715 4909 136716
rect 3371 128484 3437 128485
rect 3371 128420 3372 128484
rect 3436 128420 3437 128484
rect 3371 128419 3437 128420
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 3374 110669 3434 128419
rect 5514 115174 6134 150618
rect 6318 149837 6378 157251
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 6315 149836 6381 149837
rect 6315 149772 6316 149836
rect 6380 149772 6381 149836
rect 6315 149771 6381 149772
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3555 114068 3621 114069
rect 3555 114004 3556 114068
rect 3620 114004 3621 114068
rect 3555 114003 3621 114004
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 3558 97613 3618 114003
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 79174 6134 114618
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 8891 99652 8957 99653
rect 8891 99588 8892 99652
rect 8956 99588 8957 99652
rect 8891 99587 8957 99588
rect 8707 85236 8773 85237
rect 8707 85172 8708 85236
rect 8772 85172 8773 85236
rect 8707 85171 8773 85172
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 8710 71637 8770 85171
rect 8894 84693 8954 99587
rect 8891 84692 8957 84693
rect 8891 84628 8892 84692
rect 8956 84628 8957 84692
rect 8891 84627 8957 84628
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 8707 71636 8773 71637
rect 8707 71572 8708 71636
rect 8772 71572 8773 71636
rect 8707 71571 8773 71572
rect 8891 70820 8957 70821
rect 8891 70756 8892 70820
rect 8956 70756 8957 70820
rect 8891 70755 8957 70756
rect 8894 58581 8954 70755
rect 8891 58580 8957 58581
rect 8891 58516 8892 58580
rect 8956 58516 8957 58580
rect 8891 58515 8957 58516
rect 8891 56404 8957 56405
rect 8891 56340 8892 56404
rect 8956 56340 8957 56404
rect 8891 56339 8957 56340
rect 8894 45525 8954 56339
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 8891 45524 8957 45525
rect 8891 45460 8892 45524
rect 8956 45460 8957 45524
rect 8891 45459 8957 45460
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 8891 41988 8957 41989
rect 8891 41924 8892 41988
rect 8956 41924 8957 41988
rect 8891 41923 8957 41924
rect 8894 32469 8954 41923
rect 8891 32468 8957 32469
rect 8891 32404 8892 32468
rect 8956 32404 8957 32468
rect 8891 32403 8957 32404
rect 6315 27572 6381 27573
rect 6315 27508 6316 27572
rect 6380 27508 6381 27572
rect 6315 27507 6381 27508
rect 6318 19413 6378 27507
rect 6315 19412 6381 19413
rect 6315 19348 6316 19412
rect 6380 19348 6381 19412
rect 6315 19347 6381 19348
rect 8891 13156 8957 13157
rect 8891 13092 8892 13156
rect 8956 13092 8957 13156
rect 8891 13091 8957 13092
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 8894 6493 8954 13091
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 8891 6492 8957 6493
rect 8891 6428 8892 6492
rect 8956 6428 8957 6492
rect 8891 6427 8957 6428
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 407708 20414 416898
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 407708 24134 420618
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 407708 27854 424338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 407708 31574 428058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 407708 38414 434898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 407708 42134 438618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 407708 45854 442338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 407708 49574 410058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 407708 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 407708 60134 420618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 407708 63854 424338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 631820 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 631820 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 690600 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 690600 92414 705242
rect 95514 690600 96134 707162
rect 99234 690600 99854 709082
rect 102954 690600 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 690600 110414 704282
rect 113514 690600 114134 706202
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 690600 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 690600 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 85840 687454 86240 687486
rect 85840 687218 85922 687454
rect 86158 687218 86240 687454
rect 85840 687134 86240 687218
rect 85840 686898 85922 687134
rect 86158 686898 86240 687134
rect 85840 686866 86240 686898
rect 88440 687454 88840 687486
rect 88440 687218 88522 687454
rect 88758 687218 88840 687454
rect 88440 687134 88840 687218
rect 88440 686898 88522 687134
rect 88758 686898 88840 687134
rect 88440 686866 88840 686898
rect 95640 687454 96040 687486
rect 95640 687218 95722 687454
rect 95958 687218 96040 687454
rect 95640 687134 96040 687218
rect 95640 686898 95722 687134
rect 95958 686898 96040 687134
rect 95640 686866 96040 686898
rect 102840 687454 103240 687486
rect 102840 687218 102922 687454
rect 103158 687218 103240 687454
rect 102840 687134 103240 687218
rect 102840 686898 102922 687134
rect 103158 686898 103240 687134
rect 102840 686866 103240 686898
rect 110040 687454 110440 687486
rect 110040 687218 110122 687454
rect 110358 687218 110440 687454
rect 110040 687134 110440 687218
rect 110040 686898 110122 687134
rect 110358 686898 110440 687134
rect 110040 686866 110440 686898
rect 117240 687454 117640 687486
rect 117240 687218 117322 687454
rect 117558 687218 117640 687454
rect 117240 687134 117640 687218
rect 117240 686898 117322 687134
rect 117558 686898 117640 687134
rect 117240 686866 117640 686898
rect 119840 687454 120240 687486
rect 119840 687218 119922 687454
rect 120158 687218 120240 687454
rect 119840 687134 120240 687218
rect 119840 686898 119922 687134
rect 120158 686898 120240 687134
rect 119840 686866 120240 686898
rect 84840 669454 85240 669486
rect 84840 669218 84922 669454
rect 85158 669218 85240 669454
rect 84840 669134 85240 669218
rect 84840 668898 84922 669134
rect 85158 668898 85240 669134
rect 84840 668866 85240 668898
rect 92040 669454 92440 669486
rect 92040 669218 92122 669454
rect 92358 669218 92440 669454
rect 92040 669134 92440 669218
rect 92040 668898 92122 669134
rect 92358 668898 92440 669134
rect 92040 668866 92440 668898
rect 99240 669454 99640 669486
rect 99240 669218 99322 669454
rect 99558 669218 99640 669454
rect 99240 669134 99640 669218
rect 99240 668898 99322 669134
rect 99558 668898 99640 669134
rect 99240 668866 99640 668898
rect 106440 669454 106840 669486
rect 106440 669218 106522 669454
rect 106758 669218 106840 669454
rect 106440 669134 106840 669218
rect 106440 668898 106522 669134
rect 106758 668898 106840 669134
rect 106440 668866 106840 668898
rect 113640 669454 114040 669486
rect 113640 669218 113722 669454
rect 113958 669218 114040 669454
rect 113640 669134 114040 669218
rect 113640 668898 113722 669134
rect 113958 668898 114040 669134
rect 113640 668866 114040 668898
rect 120840 669454 121240 669486
rect 120840 669218 120922 669454
rect 121158 669218 121240 669454
rect 120840 669134 121240 669218
rect 120840 668898 120922 669134
rect 121158 668898 121240 669134
rect 120840 668866 121240 668898
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 631820 81854 658338
rect 84954 662614 85574 665600
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 631820 85574 662058
rect 91794 633454 92414 665600
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 631820 92414 632898
rect 95514 637174 96134 665600
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 631820 96134 636618
rect 99234 640894 99854 665600
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 631820 99854 640338
rect 102954 644614 103574 665600
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 631820 103574 644058
rect 109794 651454 110414 665600
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 631820 110414 650898
rect 113514 655174 114134 665600
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 631820 114134 654618
rect 117234 658894 117854 665600
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 631820 117854 658338
rect 120954 662614 121574 665600
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 631820 121574 662058
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 631820 128414 632898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 79500 615454 79820 615486
rect 79500 615218 79542 615454
rect 79778 615218 79820 615454
rect 79500 615134 79820 615218
rect 79500 614898 79542 615134
rect 79778 614898 79820 615134
rect 79500 614866 79820 614898
rect 110220 615454 110540 615486
rect 110220 615218 110262 615454
rect 110498 615218 110540 615454
rect 110220 615134 110540 615218
rect 110220 614898 110262 615134
rect 110498 614898 110540 615134
rect 110220 614866 110540 614898
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 94860 597454 95180 597486
rect 94860 597218 94902 597454
rect 95138 597218 95180 597454
rect 94860 597134 95180 597218
rect 94860 596898 94902 597134
rect 95138 596898 95180 597134
rect 94860 596866 95180 596898
rect 125580 597454 125900 597486
rect 125580 597218 125622 597454
rect 125858 597218 125900 597454
rect 125580 597134 125900 597218
rect 125580 596898 125622 597134
rect 125858 596898 125900 597134
rect 125580 596866 125900 596898
rect 79500 579454 79820 579486
rect 79500 579218 79542 579454
rect 79778 579218 79820 579454
rect 79500 579134 79820 579218
rect 79500 578898 79542 579134
rect 79778 578898 79820 579134
rect 79500 578866 79820 578898
rect 110220 579454 110540 579486
rect 110220 579218 110262 579454
rect 110498 579218 110540 579454
rect 110220 579134 110540 579218
rect 110220 578898 110262 579134
rect 110498 578898 110540 579134
rect 110220 578866 110540 578898
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 407708 67574 428058
rect 73794 543454 74414 573820
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 71083 407828 71149 407829
rect 71083 407764 71084 407828
rect 71148 407764 71149 407828
rect 71083 407763 71149 407764
rect 66115 407692 66181 407693
rect 66115 407628 66116 407692
rect 66180 407628 66181 407692
rect 66115 407627 66181 407628
rect 63539 407284 63605 407285
rect 63539 407220 63540 407284
rect 63604 407220 63605 407284
rect 63539 407219 63605 407220
rect 51027 407148 51093 407149
rect 51027 407084 51028 407148
rect 51092 407084 51093 407148
rect 51027 407083 51093 407084
rect 56179 407148 56245 407149
rect 56179 407084 56180 407148
rect 56244 407084 56245 407148
rect 56179 407083 56245 407084
rect 58571 407148 58637 407149
rect 58571 407084 58572 407148
rect 58636 407084 58637 407148
rect 58571 407083 58637 407084
rect 51030 406330 51090 407083
rect 51016 406270 51090 406330
rect 56182 406330 56242 407083
rect 58574 406330 58634 407083
rect 63542 406330 63602 407219
rect 66118 406330 66178 407627
rect 68507 407284 68573 407285
rect 68507 407220 68508 407284
rect 68572 407220 68573 407284
rect 68507 407219 68573 407220
rect 56182 406270 56244 406330
rect 48701 406196 48767 406197
rect 48701 406132 48702 406196
rect 48766 406132 48767 406196
rect 48701 406131 48767 406132
rect 48704 405620 48764 406131
rect 51016 405620 51076 406270
rect 53461 406196 53527 406197
rect 53461 406132 53462 406196
rect 53526 406132 53527 406196
rect 53461 406131 53527 406132
rect 53464 405620 53524 406131
rect 56184 405620 56244 406270
rect 58496 406270 58634 406330
rect 63528 406270 63602 406330
rect 66112 406270 66178 406330
rect 68510 406330 68570 407219
rect 71086 406330 71146 407763
rect 73794 407708 74414 434898
rect 77514 547174 78134 573820
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 407708 78134 438618
rect 81234 550894 81854 573820
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 407708 81854 442338
rect 84954 554614 85574 573820
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 407708 85574 410058
rect 91794 561454 92414 573820
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 90955 408236 91021 408237
rect 90955 408172 90956 408236
rect 91020 408172 91021 408236
rect 90955 408171 91021 408172
rect 78443 406604 78509 406605
rect 78443 406540 78444 406604
rect 78508 406540 78509 406604
rect 78443 406539 78509 406540
rect 86171 406604 86237 406605
rect 86171 406540 86172 406604
rect 86236 406540 86237 406604
rect 86171 406539 86237 406540
rect 88563 406604 88629 406605
rect 88563 406540 88564 406604
rect 88628 406540 88629 406604
rect 88563 406539 88629 406540
rect 78446 406330 78506 406539
rect 81019 406468 81085 406469
rect 81019 406404 81020 406468
rect 81084 406404 81085 406468
rect 81019 406403 81085 406404
rect 83595 406468 83661 406469
rect 83595 406404 83596 406468
rect 83660 406404 83661 406468
rect 83595 406403 83661 406404
rect 81022 406330 81082 406403
rect 68510 406270 68620 406330
rect 71086 406270 71204 406330
rect 78446 406270 78548 406330
rect 58496 405620 58556 406270
rect 61077 406196 61143 406197
rect 61077 406132 61078 406196
rect 61142 406132 61143 406196
rect 61077 406131 61143 406132
rect 61080 405620 61140 406131
rect 63528 405620 63588 406270
rect 66112 405620 66172 406270
rect 68560 405620 68620 406270
rect 71144 405620 71204 406270
rect 73589 406196 73655 406197
rect 73589 406132 73590 406196
rect 73654 406132 73655 406196
rect 73589 406131 73655 406132
rect 76173 406196 76239 406197
rect 76173 406132 76174 406196
rect 76238 406132 76239 406196
rect 76173 406131 76239 406132
rect 73592 405620 73652 406131
rect 76176 405620 76236 406131
rect 78488 405620 78548 406270
rect 80936 406270 81082 406330
rect 83598 406330 83658 406403
rect 86174 406330 86234 406539
rect 88566 406330 88626 406539
rect 83598 406270 83716 406330
rect 80936 405620 80996 406270
rect 83656 405620 83716 406270
rect 86104 406270 86234 406330
rect 88552 406270 88626 406330
rect 90958 406330 91018 408171
rect 91794 407708 92414 416898
rect 95514 565174 96134 573820
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 93531 407828 93597 407829
rect 93531 407764 93532 407828
rect 93596 407764 93597 407828
rect 93531 407763 93597 407764
rect 93534 406330 93594 407763
rect 95514 407708 96134 420618
rect 99234 568894 99854 573820
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 407708 99854 424338
rect 102954 572614 103574 573820
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 407708 103574 428058
rect 109794 543454 110414 573820
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 407708 110414 434898
rect 113514 547174 114134 573820
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 407708 114134 438618
rect 117234 550894 117854 573820
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 407708 117854 442338
rect 120954 554614 121574 573820
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 407708 121574 410058
rect 127794 561454 128414 573820
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 407708 128414 416898
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 407708 132134 420618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 407708 135854 424338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 407708 139574 428058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 139715 407964 139781 407965
rect 139715 407900 139716 407964
rect 139780 407900 139781 407964
rect 139715 407899 139781 407900
rect 101075 407692 101141 407693
rect 101075 407628 101076 407692
rect 101140 407628 101141 407692
rect 101075 407627 101141 407628
rect 98683 407148 98749 407149
rect 98683 407084 98684 407148
rect 98748 407084 98749 407148
rect 98683 407083 98749 407084
rect 95923 406604 95989 406605
rect 95923 406540 95924 406604
rect 95988 406540 95989 406604
rect 95923 406539 95989 406540
rect 90958 406270 91060 406330
rect 93534 406270 93644 406330
rect 86104 405620 86164 406270
rect 88552 405620 88612 406270
rect 91000 405620 91060 406270
rect 93584 405620 93644 406270
rect 95926 405750 95986 406539
rect 98686 405750 98746 407083
rect 101078 405750 101138 407627
rect 106043 407556 106109 407557
rect 106043 407492 106044 407556
rect 106108 407492 106109 407556
rect 106043 407491 106109 407492
rect 103651 407420 103717 407421
rect 103651 407356 103652 407420
rect 103716 407356 103717 407420
rect 103651 407355 103717 407356
rect 103654 406330 103714 407355
rect 106046 406330 106106 407491
rect 108435 407148 108501 407149
rect 108435 407084 108436 407148
rect 108500 407084 108501 407148
rect 108435 407083 108501 407084
rect 111011 407148 111077 407149
rect 111011 407084 111012 407148
rect 111076 407084 111077 407148
rect 111011 407083 111077 407084
rect 113587 407148 113653 407149
rect 113587 407084 113588 407148
rect 113652 407084 113653 407148
rect 113587 407083 113653 407084
rect 115979 407148 116045 407149
rect 115979 407084 115980 407148
rect 116044 407084 116045 407148
rect 115979 407083 116045 407084
rect 118555 407148 118621 407149
rect 118555 407084 118556 407148
rect 118620 407084 118621 407148
rect 118555 407083 118621 407084
rect 121131 407148 121197 407149
rect 121131 407084 121132 407148
rect 121196 407084 121197 407148
rect 121131 407083 121197 407084
rect 123339 407148 123405 407149
rect 123339 407084 123340 407148
rect 123404 407084 123405 407148
rect 123339 407083 123405 407084
rect 126099 407148 126165 407149
rect 126099 407084 126100 407148
rect 126164 407084 126165 407148
rect 126099 407083 126165 407084
rect 138427 407148 138493 407149
rect 138427 407084 138428 407148
rect 138492 407084 138493 407148
rect 138427 407083 138493 407084
rect 108438 406330 108498 407083
rect 111014 406330 111074 407083
rect 113590 406330 113650 407083
rect 95896 405690 95986 405750
rect 98616 405690 98746 405750
rect 101064 405690 101138 405750
rect 103512 406270 103714 406330
rect 105960 406270 106106 406330
rect 108408 406270 108498 406330
rect 110992 406270 111074 406330
rect 113576 406270 113650 406330
rect 115982 406330 116042 407083
rect 118558 406330 118618 407083
rect 121134 406330 121194 407083
rect 115982 406270 116084 406330
rect 95896 405620 95956 405690
rect 98616 405620 98676 405690
rect 101064 405620 101124 405690
rect 103512 405620 103572 406270
rect 105960 405620 106020 406270
rect 108408 405620 108468 406270
rect 110992 405620 111052 406270
rect 113576 405620 113636 406270
rect 116024 405620 116084 406270
rect 118472 406270 118618 406330
rect 121056 406270 121194 406330
rect 123342 406330 123402 407083
rect 126102 406330 126162 407083
rect 123342 406270 123428 406330
rect 118472 405620 118532 406270
rect 121056 405620 121116 406270
rect 123368 405620 123428 406270
rect 126088 406270 126162 406330
rect 138430 406330 138490 407083
rect 139718 406330 139778 407899
rect 145794 407708 146414 434898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 407708 150134 438618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 407708 153854 442338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 407708 157574 410058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 150939 407148 151005 407149
rect 150939 407084 150940 407148
rect 151004 407084 151005 407148
rect 150939 407083 151005 407084
rect 150942 406330 151002 407083
rect 138430 406270 138524 406330
rect 126088 405620 126148 406270
rect 138464 405620 138524 406270
rect 139688 406270 139778 406330
rect 150840 406270 151002 406330
rect 139688 405620 139748 406270
rect 150840 405620 150900 406270
rect 20952 399454 21300 399486
rect 20952 399218 21008 399454
rect 21244 399218 21300 399454
rect 20952 399134 21300 399218
rect 20952 398898 21008 399134
rect 21244 398898 21300 399134
rect 20952 398866 21300 398898
rect 155320 399454 155668 399486
rect 155320 399218 155376 399454
rect 155612 399218 155668 399454
rect 155320 399134 155668 399218
rect 155320 398898 155376 399134
rect 155612 398898 155668 399134
rect 155320 398866 155668 398898
rect 20272 381454 20620 381486
rect 20272 381218 20328 381454
rect 20564 381218 20620 381454
rect 20272 381134 20620 381218
rect 20272 380898 20328 381134
rect 20564 380898 20620 381134
rect 20272 380866 20620 380898
rect 156000 381454 156348 381486
rect 156000 381218 156056 381454
rect 156292 381218 156348 381454
rect 156000 381134 156348 381218
rect 156000 380898 156056 381134
rect 156292 380898 156348 381134
rect 156000 380866 156348 380898
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 20952 363454 21300 363486
rect 20952 363218 21008 363454
rect 21244 363218 21300 363454
rect 20952 363134 21300 363218
rect 20952 362898 21008 363134
rect 21244 362898 21300 363134
rect 20952 362866 21300 362898
rect 155320 363454 155668 363486
rect 155320 363218 155376 363454
rect 155612 363218 155668 363454
rect 155320 363134 155668 363218
rect 155320 362898 155376 363134
rect 155612 362898 155668 363134
rect 155320 362866 155668 362898
rect 20272 345454 20620 345486
rect 20272 345218 20328 345454
rect 20564 345218 20620 345454
rect 20272 345134 20620 345218
rect 20272 344898 20328 345134
rect 20564 344898 20620 345134
rect 20272 344866 20620 344898
rect 156000 345454 156348 345486
rect 156000 345218 156056 345454
rect 156292 345218 156348 345454
rect 156000 345134 156348 345218
rect 156000 344898 156056 345134
rect 156292 344898 156348 345134
rect 156000 344866 156348 344898
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 20952 327454 21300 327486
rect 20952 327218 21008 327454
rect 21244 327218 21300 327454
rect 20952 327134 21300 327218
rect 20952 326898 21008 327134
rect 21244 326898 21300 327134
rect 20952 326866 21300 326898
rect 155320 327454 155668 327486
rect 155320 327218 155376 327454
rect 155612 327218 155668 327454
rect 155320 327134 155668 327218
rect 155320 326898 155376 327134
rect 155612 326898 155668 327134
rect 155320 326866 155668 326898
rect 36056 322010 36116 322506
rect 37144 322010 37204 322506
rect 36056 321950 36186 322010
rect 19011 321468 19077 321469
rect 19011 321404 19012 321468
rect 19076 321404 19077 321468
rect 19011 321403 19077 321404
rect 18827 319836 18893 319837
rect 18827 319772 18828 319836
rect 18892 319772 18893 319836
rect 18827 319771 18893 319772
rect 18643 319564 18709 319565
rect 18643 319500 18644 319564
rect 18708 319500 18709 319564
rect 18643 319499 18709 319500
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 18459 287740 18525 287741
rect 18459 287676 18460 287740
rect 18524 287676 18525 287740
rect 18459 287675 18525 287676
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 18462 200293 18522 287675
rect 18646 200701 18706 319499
rect 18643 200700 18709 200701
rect 18643 200636 18644 200700
rect 18708 200636 18709 200700
rect 18643 200635 18709 200636
rect 18830 200429 18890 319771
rect 19014 201109 19074 321403
rect 19195 321332 19261 321333
rect 19195 321268 19196 321332
rect 19260 321268 19261 321332
rect 19195 321267 19261 321268
rect 19011 201108 19077 201109
rect 19011 201044 19012 201108
rect 19076 201044 19077 201108
rect 19011 201043 19077 201044
rect 19198 200973 19258 321267
rect 19379 320652 19445 320653
rect 19379 320588 19380 320652
rect 19444 320588 19445 320652
rect 19379 320587 19445 320588
rect 19382 316029 19442 320587
rect 20667 320516 20733 320517
rect 20667 320452 20668 320516
rect 20732 320452 20733 320516
rect 20667 320451 20733 320452
rect 19563 319428 19629 319429
rect 19563 319364 19564 319428
rect 19628 319364 19629 319428
rect 19563 319363 19629 319364
rect 19566 316301 19626 319363
rect 19563 316300 19629 316301
rect 19563 316236 19564 316300
rect 19628 316236 19629 316300
rect 19563 316235 19629 316236
rect 19563 316164 19629 316165
rect 19563 316100 19564 316164
rect 19628 316100 19629 316164
rect 19563 316099 19629 316100
rect 19379 316028 19445 316029
rect 19379 315964 19380 316028
rect 19444 315964 19445 316028
rect 19379 315963 19445 315964
rect 19379 315892 19445 315893
rect 19379 315828 19380 315892
rect 19444 315828 19445 315892
rect 19379 315827 19445 315828
rect 19382 306645 19442 315827
rect 19379 306644 19445 306645
rect 19379 306580 19380 306644
rect 19444 306580 19445 306644
rect 19379 306579 19445 306580
rect 19379 306508 19445 306509
rect 19379 306444 19380 306508
rect 19444 306444 19445 306508
rect 19379 306443 19445 306444
rect 19382 306373 19442 306443
rect 19379 306372 19445 306373
rect 19379 306308 19380 306372
rect 19444 306308 19445 306372
rect 19379 306307 19445 306308
rect 19379 306236 19445 306237
rect 19379 306172 19380 306236
rect 19444 306172 19445 306236
rect 19379 306171 19445 306172
rect 19382 296989 19442 306171
rect 19379 296988 19445 296989
rect 19379 296924 19380 296988
rect 19444 296924 19445 296988
rect 19379 296923 19445 296924
rect 19379 296852 19445 296853
rect 19379 296788 19380 296852
rect 19444 296788 19445 296852
rect 19379 296787 19445 296788
rect 19382 296717 19442 296787
rect 19379 296716 19445 296717
rect 19379 296652 19380 296716
rect 19444 296652 19445 296716
rect 19379 296651 19445 296652
rect 19379 296580 19445 296581
rect 19379 296516 19380 296580
rect 19444 296516 19445 296580
rect 19379 296515 19445 296516
rect 19382 288965 19442 296515
rect 19379 288964 19445 288965
rect 19379 288900 19380 288964
rect 19444 288900 19445 288964
rect 19379 288899 19445 288900
rect 19379 288556 19445 288557
rect 19379 288492 19380 288556
rect 19444 288492 19445 288556
rect 19379 288491 19445 288492
rect 19195 200972 19261 200973
rect 19195 200908 19196 200972
rect 19260 200908 19261 200972
rect 19195 200907 19261 200908
rect 19382 200565 19442 288491
rect 19566 200837 19626 316099
rect 19794 309454 20414 320400
rect 20670 316050 20730 320451
rect 20670 315990 20914 316050
rect 20667 315892 20733 315893
rect 20667 315828 20668 315892
rect 20732 315828 20733 315892
rect 20667 315827 20733 315828
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 289308 20414 308898
rect 20670 296853 20730 315827
rect 20854 306509 20914 315990
rect 23514 313174 24134 320400
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 20851 306508 20917 306509
rect 20851 306444 20852 306508
rect 20916 306444 20917 306508
rect 20851 306443 20917 306444
rect 20851 306372 20917 306373
rect 20851 306308 20852 306372
rect 20916 306308 20917 306372
rect 20851 306307 20917 306308
rect 20667 296852 20733 296853
rect 20667 296788 20668 296852
rect 20732 296788 20733 296852
rect 20667 296787 20733 296788
rect 20667 296580 20733 296581
rect 20667 296516 20668 296580
rect 20732 296516 20733 296580
rect 20667 296515 20733 296516
rect 19747 288964 19813 288965
rect 19747 288900 19748 288964
rect 19812 288900 19813 288964
rect 19747 288899 19813 288900
rect 19750 202877 19810 288899
rect 20670 288690 20730 296515
rect 19934 288630 20730 288690
rect 19934 203690 19994 288630
rect 20854 288557 20914 306307
rect 23514 289308 24134 312618
rect 27234 316894 27854 320400
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 289308 27854 316338
rect 30954 301674 31574 320400
rect 36126 319973 36186 321950
rect 37046 321950 37204 322010
rect 38232 322010 38292 322506
rect 39592 322010 39652 322506
rect 40544 322010 40604 322506
rect 38232 321950 38578 322010
rect 39592 321950 39682 322010
rect 36123 319972 36189 319973
rect 36123 319908 36124 319972
rect 36188 319908 36189 319972
rect 36123 319907 36189 319908
rect 37046 319157 37106 321950
rect 37043 319156 37109 319157
rect 37043 319092 37044 319156
rect 37108 319092 37109 319156
rect 37043 319091 37109 319092
rect 30954 301438 30986 301674
rect 31222 301438 31306 301674
rect 31542 301438 31574 301674
rect 30954 301354 31574 301438
rect 30954 301118 30986 301354
rect 31222 301118 31306 301354
rect 31542 301118 31574 301354
rect 30954 289308 31574 301118
rect 37794 291454 38414 320400
rect 38518 319157 38578 321950
rect 39622 319973 39682 321950
rect 40542 321950 40604 322010
rect 41768 322010 41828 322506
rect 43128 322010 43188 322506
rect 41768 321950 42442 322010
rect 39619 319972 39685 319973
rect 39619 319908 39620 319972
rect 39684 319908 39685 319972
rect 39619 319907 39685 319908
rect 40542 319293 40602 321950
rect 40539 319292 40605 319293
rect 40539 319228 40540 319292
rect 40604 319228 40605 319292
rect 40539 319227 40605 319228
rect 38515 319156 38581 319157
rect 38515 319092 38516 319156
rect 38580 319092 38581 319156
rect 38515 319091 38581 319092
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 289308 38414 290898
rect 41514 295174 42134 320400
rect 42382 319293 42442 321950
rect 43118 321950 43188 322010
rect 44216 322010 44276 322506
rect 45440 322010 45500 322506
rect 46528 322010 46588 322506
rect 47616 322010 47676 322506
rect 48704 322010 48764 322506
rect 44216 321950 44282 322010
rect 43118 320245 43178 321950
rect 43115 320244 43181 320245
rect 43115 320180 43116 320244
rect 43180 320180 43181 320244
rect 43115 320179 43181 320180
rect 44222 320109 44282 321950
rect 44958 321950 45500 322010
rect 46430 321950 46588 322010
rect 47534 321950 47676 322010
rect 48638 321950 48764 322010
rect 50064 322010 50124 322506
rect 51288 322010 51348 322506
rect 52376 322010 52436 322506
rect 53464 322010 53524 322506
rect 54552 322010 54612 322506
rect 55912 322010 55972 322506
rect 57000 322010 57060 322506
rect 50064 321950 50170 322010
rect 44958 320109 45018 321950
rect 44219 320108 44285 320109
rect 44219 320044 44220 320108
rect 44284 320044 44285 320108
rect 44219 320043 44285 320044
rect 44955 320108 45021 320109
rect 44955 320044 44956 320108
rect 45020 320044 45021 320108
rect 44955 320043 45021 320044
rect 42379 319292 42445 319293
rect 42379 319228 42380 319292
rect 42444 319228 42445 319292
rect 42379 319227 42445 319228
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 289308 42134 294618
rect 45234 298894 45854 320400
rect 46430 319157 46490 321950
rect 47534 319429 47594 321950
rect 48638 319565 48698 321950
rect 48635 319564 48701 319565
rect 48635 319500 48636 319564
rect 48700 319500 48701 319564
rect 48635 319499 48701 319500
rect 47531 319428 47597 319429
rect 47531 319364 47532 319428
rect 47596 319364 47597 319428
rect 47531 319363 47597 319364
rect 46427 319156 46493 319157
rect 46427 319092 46428 319156
rect 46492 319092 46493 319156
rect 46427 319091 46493 319092
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 289308 45854 298338
rect 48954 302614 49574 320400
rect 50110 320109 50170 321950
rect 51214 321950 51348 322010
rect 52318 321950 52436 322010
rect 53422 321950 53524 322010
rect 54526 321950 54612 322010
rect 55630 321950 55972 322010
rect 56918 321950 57060 322010
rect 58088 322010 58148 322506
rect 59448 322010 59508 322506
rect 60672 322010 60732 322506
rect 61760 322010 61820 322506
rect 62848 322010 62908 322506
rect 63936 322010 63996 322506
rect 58088 321950 58266 322010
rect 51214 320109 51274 321950
rect 52318 320109 52378 321950
rect 53422 320109 53482 321950
rect 54526 321197 54586 321950
rect 54523 321196 54589 321197
rect 54523 321132 54524 321196
rect 54588 321132 54589 321196
rect 54523 321131 54589 321132
rect 50107 320108 50173 320109
rect 50107 320044 50108 320108
rect 50172 320044 50173 320108
rect 50107 320043 50173 320044
rect 51211 320108 51277 320109
rect 51211 320044 51212 320108
rect 51276 320044 51277 320108
rect 51211 320043 51277 320044
rect 52315 320108 52381 320109
rect 52315 320044 52316 320108
rect 52380 320044 52381 320108
rect 52315 320043 52381 320044
rect 53419 320108 53485 320109
rect 53419 320044 53420 320108
rect 53484 320044 53485 320108
rect 53419 320043 53485 320044
rect 55630 319701 55690 321950
rect 56918 321333 56978 321950
rect 58206 321469 58266 321950
rect 59310 321950 59508 322010
rect 60598 321950 60732 322010
rect 61702 321950 61820 322010
rect 62806 321950 62908 322010
rect 63910 321950 63996 322010
rect 65296 322010 65356 322506
rect 66384 322010 66444 322506
rect 67608 322010 67668 322506
rect 68696 322010 68756 322506
rect 65296 321950 65442 322010
rect 66384 321950 66546 322010
rect 58203 321468 58269 321469
rect 58203 321404 58204 321468
rect 58268 321404 58269 321468
rect 58203 321403 58269 321404
rect 56915 321332 56981 321333
rect 56915 321268 56916 321332
rect 56980 321268 56981 321332
rect 56915 321267 56981 321268
rect 55627 319700 55693 319701
rect 55627 319636 55628 319700
rect 55692 319636 55693 319700
rect 55627 319635 55693 319636
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48635 291140 48701 291141
rect 48635 291076 48636 291140
rect 48700 291076 48701 291140
rect 48635 291075 48701 291076
rect 20851 288556 20917 288557
rect 20851 288492 20852 288556
rect 20916 288492 20917 288556
rect 20851 288491 20917 288492
rect 48638 288010 48698 291075
rect 48954 289308 49574 302058
rect 55794 309454 56414 320400
rect 59310 320109 59370 321950
rect 59307 320108 59373 320109
rect 59307 320044 59308 320108
rect 59372 320044 59373 320108
rect 59307 320043 59373 320044
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 51027 291140 51093 291141
rect 51027 291076 51028 291140
rect 51092 291076 51093 291140
rect 51027 291075 51093 291076
rect 53419 291140 53485 291141
rect 53419 291076 53420 291140
rect 53484 291076 53485 291140
rect 53419 291075 53485 291076
rect 51030 288010 51090 291075
rect 48638 287950 48764 288010
rect 48704 287300 48764 287950
rect 51016 287950 51090 288010
rect 53422 288010 53482 291075
rect 55794 289308 56414 308898
rect 59514 313174 60134 320400
rect 60598 319973 60658 321950
rect 61702 320653 61762 321950
rect 62806 321605 62866 321950
rect 63910 321605 63970 321950
rect 62803 321604 62869 321605
rect 62803 321540 62804 321604
rect 62868 321540 62869 321604
rect 62803 321539 62869 321540
rect 63907 321604 63973 321605
rect 63907 321540 63908 321604
rect 63972 321540 63973 321604
rect 63907 321539 63973 321540
rect 61699 320652 61765 320653
rect 61699 320588 61700 320652
rect 61764 320588 61765 320652
rect 61699 320587 61765 320588
rect 60595 319972 60661 319973
rect 60595 319908 60596 319972
rect 60660 319908 60661 319972
rect 60595 319907 60661 319908
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 56547 291140 56613 291141
rect 56547 291076 56548 291140
rect 56612 291076 56613 291140
rect 56547 291075 56613 291076
rect 58571 291140 58637 291141
rect 58571 291076 58572 291140
rect 58636 291076 58637 291140
rect 58571 291075 58637 291076
rect 56550 288010 56610 291075
rect 58574 288010 58634 291075
rect 59514 289308 60134 312618
rect 63234 316894 63854 320400
rect 65382 320109 65442 321950
rect 66486 321741 66546 321950
rect 67590 321950 67668 322010
rect 68694 321950 68756 322010
rect 69784 322010 69844 322506
rect 71144 322010 71204 322506
rect 72232 322010 72292 322506
rect 73320 322010 73380 322506
rect 74408 322010 74468 322506
rect 75768 322010 75828 322506
rect 76992 322010 77052 322506
rect 69784 321950 69858 322010
rect 66483 321740 66549 321741
rect 66483 321676 66484 321740
rect 66548 321676 66549 321740
rect 66483 321675 66549 321676
rect 65379 320108 65445 320109
rect 65379 320044 65380 320108
rect 65444 320044 65445 320108
rect 65379 320043 65445 320044
rect 66486 319973 66546 321675
rect 67590 321605 67650 321950
rect 68694 321877 68754 321950
rect 68691 321876 68757 321877
rect 68691 321812 68692 321876
rect 68756 321812 68757 321876
rect 68691 321811 68757 321812
rect 67587 321604 67653 321605
rect 67587 321540 67588 321604
rect 67652 321540 67653 321604
rect 67587 321539 67653 321540
rect 66483 319972 66549 319973
rect 66483 319908 66484 319972
rect 66548 319908 66549 319972
rect 66483 319907 66549 319908
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 61147 291140 61213 291141
rect 61147 291076 61148 291140
rect 61212 291076 61213 291140
rect 61147 291075 61213 291076
rect 61150 288010 61210 291075
rect 63234 289308 63854 316338
rect 66954 301674 67574 320400
rect 68694 320109 68754 321811
rect 68691 320108 68757 320109
rect 68691 320044 68692 320108
rect 68756 320044 68757 320108
rect 68691 320043 68757 320044
rect 69798 319293 69858 321950
rect 71086 321950 71204 322010
rect 72190 321950 72292 322010
rect 73294 321950 73380 322010
rect 74398 321950 74468 322010
rect 75686 321950 75828 322010
rect 76974 321950 77052 322010
rect 78080 322010 78140 322506
rect 79168 322010 79228 322506
rect 143224 322010 143284 322506
rect 143360 322013 143420 322506
rect 78080 321950 78322 322010
rect 79168 321950 79242 322010
rect 71086 320109 71146 321950
rect 72190 320109 72250 321950
rect 73294 320109 73354 321950
rect 74398 320650 74458 321950
rect 74398 320590 74642 320650
rect 74582 320517 74642 320590
rect 74579 320516 74645 320517
rect 74579 320452 74580 320516
rect 74644 320452 74645 320516
rect 74579 320451 74645 320452
rect 71083 320108 71149 320109
rect 71083 320044 71084 320108
rect 71148 320044 71149 320108
rect 71083 320043 71149 320044
rect 72187 320108 72253 320109
rect 72187 320044 72188 320108
rect 72252 320044 72253 320108
rect 72187 320043 72253 320044
rect 73291 320108 73357 320109
rect 73291 320044 73292 320108
rect 73356 320044 73357 320108
rect 73291 320043 73357 320044
rect 69795 319292 69861 319293
rect 69795 319228 69796 319292
rect 69860 319228 69861 319292
rect 69795 319227 69861 319228
rect 66954 301438 66986 301674
rect 67222 301438 67306 301674
rect 67542 301438 67574 301674
rect 66954 301354 67574 301438
rect 66954 301118 66986 301354
rect 67222 301118 67306 301354
rect 67542 301118 67574 301354
rect 64091 291140 64157 291141
rect 64091 291076 64092 291140
rect 64156 291076 64157 291140
rect 64091 291075 64157 291076
rect 64094 288010 64154 291075
rect 64827 290732 64893 290733
rect 64827 290730 64828 290732
rect 53422 287950 53524 288010
rect 51016 287300 51076 287950
rect 53464 287300 53524 287950
rect 56184 287950 56610 288010
rect 58496 287950 58634 288010
rect 61080 287950 61210 288010
rect 63528 287950 64154 288010
rect 64646 290670 64828 290730
rect 64646 288010 64706 290670
rect 64827 290668 64828 290670
rect 64892 290668 64893 290732
rect 64827 290667 64893 290668
rect 66954 289308 67574 301118
rect 73794 291454 74414 320400
rect 75686 320109 75746 321950
rect 75683 320108 75749 320109
rect 75683 320044 75684 320108
rect 75748 320044 75749 320108
rect 75683 320043 75749 320044
rect 76974 319293 77034 321950
rect 76971 319292 77037 319293
rect 76971 319228 76972 319292
rect 77036 319228 77037 319292
rect 76971 319227 77037 319228
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 68507 291140 68573 291141
rect 68507 291076 68508 291140
rect 68572 291076 68573 291140
rect 68507 291075 68573 291076
rect 71083 291140 71149 291141
rect 71083 291076 71084 291140
rect 71148 291076 71149 291140
rect 71083 291075 71149 291076
rect 73794 291134 74414 291218
rect 77514 295174 78134 320400
rect 78262 319701 78322 321950
rect 79182 320109 79242 321950
rect 143214 321950 143284 322010
rect 143357 322012 143423 322013
rect 143214 320517 143274 321950
rect 143357 321948 143358 322012
rect 143422 321948 143423 322012
rect 143357 321947 143423 321948
rect 143211 320516 143277 320517
rect 143211 320452 143212 320516
rect 143276 320452 143277 320516
rect 143211 320451 143277 320452
rect 79179 320108 79245 320109
rect 79179 320044 79180 320108
rect 79244 320044 79245 320108
rect 79179 320043 79245 320044
rect 78259 319700 78325 319701
rect 78259 319636 78260 319700
rect 78324 319636 78325 319700
rect 78259 319635 78325 319636
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 68510 288010 68570 291075
rect 71086 288010 71146 291075
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 76235 291140 76301 291141
rect 76235 291076 76236 291140
rect 76300 291076 76301 291140
rect 76235 291075 76301 291076
rect 73475 290324 73541 290325
rect 73475 290260 73476 290324
rect 73540 290260 73541 290324
rect 73475 290259 73541 290260
rect 73478 288010 73538 290259
rect 73794 289308 74414 290898
rect 76238 288010 76298 291075
rect 77514 289308 78134 294618
rect 81234 298894 81854 320400
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 78443 291140 78509 291141
rect 78443 291076 78444 291140
rect 78508 291076 78509 291140
rect 78443 291075 78509 291076
rect 81019 291140 81085 291141
rect 81019 291076 81020 291140
rect 81084 291076 81085 291140
rect 81019 291075 81085 291076
rect 64646 287950 66172 288010
rect 68510 287950 68620 288010
rect 71086 287950 71204 288010
rect 73478 287950 73652 288010
rect 56184 287300 56244 287950
rect 58496 287300 58556 287950
rect 61080 287300 61140 287950
rect 63528 287300 63588 287950
rect 66112 287300 66172 287950
rect 68560 287300 68620 287950
rect 71144 287300 71204 287950
rect 73592 287300 73652 287950
rect 76176 287950 76298 288010
rect 78446 288010 78506 291075
rect 81022 288010 81082 291075
rect 81234 289308 81854 298338
rect 84954 302614 85574 320400
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 83595 291140 83661 291141
rect 83595 291076 83596 291140
rect 83660 291076 83661 291140
rect 83595 291075 83661 291076
rect 78446 287950 78548 288010
rect 76176 287300 76236 287950
rect 78488 287300 78548 287950
rect 80936 287950 81082 288010
rect 83598 288010 83658 291075
rect 84954 289308 85574 302058
rect 91794 309454 92414 320400
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 86171 291140 86237 291141
rect 86171 291076 86172 291140
rect 86236 291076 86237 291140
rect 86171 291075 86237 291076
rect 88563 291140 88629 291141
rect 88563 291076 88564 291140
rect 88628 291076 88629 291140
rect 88563 291075 88629 291076
rect 90955 291140 91021 291141
rect 90955 291076 90956 291140
rect 91020 291076 91021 291140
rect 90955 291075 91021 291076
rect 86174 288010 86234 291075
rect 88566 288010 88626 291075
rect 83598 287950 83716 288010
rect 80936 287300 80996 287950
rect 83656 287300 83716 287950
rect 86104 287950 86234 288010
rect 88552 287950 88626 288010
rect 90958 288010 91018 291075
rect 91794 289308 92414 308898
rect 95514 313174 96134 320400
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 93531 291140 93597 291141
rect 93531 291076 93532 291140
rect 93596 291076 93597 291140
rect 93531 291075 93597 291076
rect 93534 288010 93594 291075
rect 95514 289308 96134 312618
rect 99234 316894 99854 320400
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 98683 291140 98749 291141
rect 98683 291076 98684 291140
rect 98748 291076 98749 291140
rect 98683 291075 98749 291076
rect 96291 290188 96357 290189
rect 96291 290124 96292 290188
rect 96356 290124 96357 290188
rect 96291 290123 96357 290124
rect 96294 288010 96354 290123
rect 98686 288010 98746 291075
rect 99234 289308 99854 316338
rect 102954 301674 103574 320400
rect 102954 301438 102986 301674
rect 103222 301438 103306 301674
rect 103542 301438 103574 301674
rect 102954 301354 103574 301438
rect 102954 301118 102986 301354
rect 103222 301118 103306 301354
rect 103542 301118 103574 301354
rect 101075 291004 101141 291005
rect 101075 290940 101076 291004
rect 101140 290940 101141 291004
rect 101075 290939 101141 290940
rect 101078 288010 101138 290939
rect 102954 289308 103574 301118
rect 109794 291454 110414 320400
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 106043 291140 106109 291141
rect 106043 291076 106044 291140
rect 106108 291076 106109 291140
rect 106043 291075 106109 291076
rect 109794 291134 110414 291218
rect 103835 290732 103901 290733
rect 103835 290668 103836 290732
rect 103900 290668 103901 290732
rect 103835 290667 103901 290668
rect 103838 288010 103898 290667
rect 106046 288010 106106 291075
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 113514 295174 114134 320400
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113219 291004 113285 291005
rect 113219 290940 113220 291004
rect 113284 290940 113285 291004
rect 113219 290939 113285 290940
rect 108435 290052 108501 290053
rect 108435 289988 108436 290052
rect 108500 289988 108501 290052
rect 108435 289987 108501 289988
rect 108438 288010 108498 289987
rect 109794 289308 110414 290898
rect 111011 290868 111077 290869
rect 111011 290804 111012 290868
rect 111076 290804 111077 290868
rect 111011 290803 111077 290804
rect 111014 288010 111074 290803
rect 90958 287950 91060 288010
rect 93534 287950 93644 288010
rect 86104 287300 86164 287950
rect 88552 287300 88612 287950
rect 91000 287300 91060 287950
rect 93584 287300 93644 287950
rect 95896 287950 96354 288010
rect 98616 287950 98746 288010
rect 101064 287950 101138 288010
rect 103512 287950 103898 288010
rect 105960 287950 106106 288010
rect 108408 287950 108498 288010
rect 110992 287950 111074 288010
rect 113222 288010 113282 290939
rect 113514 289308 114134 294618
rect 117234 298894 117854 320400
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 115979 291140 116045 291141
rect 115979 291076 115980 291140
rect 116044 291076 116045 291140
rect 115979 291075 116045 291076
rect 115982 288010 116042 291075
rect 117234 289308 117854 298338
rect 120954 302614 121574 320400
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 118555 290732 118621 290733
rect 118555 290668 118556 290732
rect 118620 290668 118621 290732
rect 118555 290667 118621 290668
rect 118558 288010 118618 290667
rect 120763 290324 120829 290325
rect 120763 290260 120764 290324
rect 120828 290260 120829 290324
rect 120763 290259 120829 290260
rect 113222 287950 113636 288010
rect 115982 287950 116084 288010
rect 95896 287300 95956 287950
rect 98616 287300 98676 287950
rect 101064 287300 101124 287950
rect 103512 287300 103572 287950
rect 105960 287300 106020 287950
rect 108408 287300 108468 287950
rect 110992 287300 111052 287950
rect 113576 287300 113636 287950
rect 116024 287300 116084 287950
rect 118472 287950 118618 288010
rect 120766 288010 120826 290259
rect 120954 289308 121574 302058
rect 127794 309454 128414 320400
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 126099 290460 126165 290461
rect 126099 290396 126100 290460
rect 126164 290396 126165 290460
rect 126099 290395 126165 290396
rect 122787 290052 122853 290053
rect 122787 290050 122788 290052
rect 122606 289990 122788 290050
rect 122606 288010 122666 289990
rect 122787 289988 122788 289990
rect 122852 289988 122853 290052
rect 122787 289987 122853 289988
rect 126102 288010 126162 290395
rect 127794 289308 128414 308898
rect 131514 313174 132134 320400
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 289308 132134 312618
rect 135234 316894 135854 320400
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 289308 135854 316338
rect 138954 301674 139574 320400
rect 138954 301438 138986 301674
rect 139222 301438 139306 301674
rect 139542 301438 139574 301674
rect 138954 301354 139574 301438
rect 138954 301118 138986 301354
rect 139222 301118 139306 301354
rect 139542 301118 139574 301354
rect 138427 290460 138493 290461
rect 138427 290396 138428 290460
rect 138492 290396 138493 290460
rect 138427 290395 138493 290396
rect 120766 287950 121116 288010
rect 122606 287950 123428 288010
rect 118472 287300 118532 287950
rect 121056 287300 121116 287950
rect 123368 287300 123428 287950
rect 126088 287950 126162 288010
rect 138430 288010 138490 290395
rect 138954 289308 139574 301118
rect 145794 291454 146414 320400
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 139715 290868 139781 290869
rect 139715 290804 139716 290868
rect 139780 290804 139781 290868
rect 139715 290803 139781 290804
rect 139718 288010 139778 290803
rect 145794 289308 146414 290898
rect 149514 295174 150134 320400
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 289308 150134 294618
rect 153234 298894 153854 320400
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 289308 153854 298338
rect 156954 302614 157574 320400
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 289308 157574 302058
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 138430 287950 138524 288010
rect 126088 287300 126148 287950
rect 138464 287300 138524 287950
rect 139688 287950 139778 288010
rect 139688 287300 139748 287950
rect 150837 287468 150903 287469
rect 150837 287404 150838 287468
rect 150902 287404 150903 287468
rect 150837 287403 150903 287404
rect 150840 287300 150900 287403
rect 20272 273454 20620 273486
rect 20272 273218 20328 273454
rect 20564 273218 20620 273454
rect 20272 273134 20620 273218
rect 20272 272898 20328 273134
rect 20564 272898 20620 273134
rect 20272 272866 20620 272898
rect 156000 273454 156348 273486
rect 156000 273218 156056 273454
rect 156292 273218 156348 273454
rect 156000 273134 156348 273218
rect 156000 272898 156056 273134
rect 156292 272898 156348 273134
rect 156000 272866 156348 272898
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 20952 255454 21300 255486
rect 20952 255218 21008 255454
rect 21244 255218 21300 255454
rect 20952 255134 21300 255218
rect 20952 254898 21008 255134
rect 21244 254898 21300 255134
rect 20952 254866 21300 254898
rect 155320 255454 155668 255486
rect 155320 255218 155376 255454
rect 155612 255218 155668 255454
rect 155320 255134 155668 255218
rect 155320 254898 155376 255134
rect 155612 254898 155668 255134
rect 155320 254866 155668 254898
rect 20272 237454 20620 237486
rect 20272 237218 20328 237454
rect 20564 237218 20620 237454
rect 20272 237134 20620 237218
rect 20272 236898 20328 237134
rect 20564 236898 20620 237134
rect 20272 236866 20620 236898
rect 156000 237454 156348 237486
rect 156000 237218 156056 237454
rect 156292 237218 156348 237454
rect 156000 237134 156348 237218
rect 156000 236898 156056 237134
rect 156292 236898 156348 237134
rect 156000 236866 156348 236898
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 20952 219454 21300 219486
rect 20952 219218 21008 219454
rect 21244 219218 21300 219454
rect 20952 219134 21300 219218
rect 20952 218898 21008 219134
rect 21244 218898 21300 219134
rect 20952 218866 21300 218898
rect 155320 219454 155668 219486
rect 155320 219218 155376 219454
rect 155612 219218 155668 219454
rect 155320 219134 155668 219218
rect 155320 218898 155376 219134
rect 155612 218898 155668 219134
rect 155320 218866 155668 218898
rect 36056 203690 36116 204000
rect 37144 203690 37204 204000
rect 19934 203630 20730 203690
rect 19747 202876 19813 202877
rect 19747 202812 19748 202876
rect 19812 202812 19813 202876
rect 19747 202811 19813 202812
rect 19794 201454 20414 202000
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 20670 201245 20730 203630
rect 35942 203630 36116 203690
rect 37046 203630 37204 203690
rect 38232 203690 38292 204000
rect 39592 203690 39652 204000
rect 40544 203690 40604 204000
rect 41768 203690 41828 204000
rect 43128 203690 43188 204000
rect 38232 203630 38578 203690
rect 39592 203630 39682 203690
rect 19794 201134 20414 201218
rect 20667 201244 20733 201245
rect 20667 201180 20668 201244
rect 20732 201180 20733 201244
rect 20667 201179 20733 201180
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19563 200836 19629 200837
rect 19563 200772 19564 200836
rect 19628 200772 19629 200836
rect 19563 200771 19629 200772
rect 19379 200564 19445 200565
rect 19379 200500 19380 200564
rect 19444 200500 19445 200564
rect 19379 200499 19445 200500
rect 18827 200428 18893 200429
rect 18827 200364 18828 200428
rect 18892 200364 18893 200428
rect 18827 200363 18893 200364
rect 18459 200292 18525 200293
rect 18459 200228 18460 200292
rect 18524 200228 18525 200292
rect 18459 200227 18525 200228
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 169174 24134 202000
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 172894 27854 202000
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 176614 31574 202000
rect 35942 201381 36002 203630
rect 37046 201381 37106 203630
rect 35939 201380 36005 201381
rect 35939 201316 35940 201380
rect 36004 201316 36005 201380
rect 35939 201315 36005 201316
rect 37043 201380 37109 201381
rect 37043 201316 37044 201380
rect 37108 201316 37109 201380
rect 37043 201315 37109 201316
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 183454 38414 202000
rect 38518 201381 38578 203630
rect 39622 201381 39682 203630
rect 40542 203630 40604 203690
rect 41646 203630 41828 203690
rect 43118 203630 43188 203690
rect 44216 203690 44276 204000
rect 45440 203690 45500 204000
rect 46528 203690 46588 204000
rect 47616 203690 47676 204000
rect 48704 203690 48764 204000
rect 44216 203630 44282 203690
rect 40542 201381 40602 203630
rect 41646 202197 41706 203630
rect 41643 202196 41709 202197
rect 41643 202132 41644 202196
rect 41708 202132 41709 202196
rect 41643 202131 41709 202132
rect 38515 201380 38581 201381
rect 38515 201316 38516 201380
rect 38580 201316 38581 201380
rect 38515 201315 38581 201316
rect 39619 201380 39685 201381
rect 39619 201316 39620 201380
rect 39684 201316 39685 201380
rect 39619 201315 39685 201316
rect 40539 201380 40605 201381
rect 40539 201316 40540 201380
rect 40604 201316 40605 201380
rect 40539 201315 40605 201316
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 187174 42134 202000
rect 43118 200429 43178 203630
rect 44222 201381 44282 203630
rect 44958 203630 45500 203690
rect 46430 203630 46588 203690
rect 47534 203630 47676 203690
rect 48638 203630 48764 203690
rect 50064 203690 50124 204000
rect 51288 203690 51348 204000
rect 52376 203690 52436 204000
rect 53464 203690 53524 204000
rect 54552 203690 54612 204000
rect 55912 203690 55972 204000
rect 57000 203690 57060 204000
rect 58088 203690 58148 204000
rect 59448 203690 59508 204000
rect 60672 203690 60732 204000
rect 61760 203690 61820 204000
rect 62848 203690 62908 204000
rect 50064 203630 50170 203690
rect 44958 201381 45018 203630
rect 44219 201380 44285 201381
rect 44219 201316 44220 201380
rect 44284 201316 44285 201380
rect 44219 201315 44285 201316
rect 44955 201380 45021 201381
rect 44955 201316 44956 201380
rect 45020 201316 45021 201380
rect 44955 201315 45021 201316
rect 43115 200428 43181 200429
rect 43115 200364 43116 200428
rect 43180 200364 43181 200428
rect 43115 200363 43181 200364
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 190894 45854 202000
rect 46430 200293 46490 203630
rect 47534 202877 47594 203630
rect 47531 202876 47597 202877
rect 47531 202812 47532 202876
rect 47596 202812 47597 202876
rect 47531 202811 47597 202812
rect 48638 200701 48698 203630
rect 48635 200700 48701 200701
rect 48635 200636 48636 200700
rect 48700 200636 48701 200700
rect 48635 200635 48701 200636
rect 46427 200292 46493 200293
rect 46427 200228 46428 200292
rect 46492 200228 46493 200292
rect 46427 200227 46493 200228
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 194614 49574 202000
rect 50110 200837 50170 203630
rect 51214 203630 51348 203690
rect 52318 203630 52436 203690
rect 53422 203630 53524 203690
rect 54526 203630 54612 203690
rect 55630 203630 55972 203690
rect 56918 203630 57060 203690
rect 58022 203630 58148 203690
rect 59310 203630 59508 203690
rect 60598 203630 60732 203690
rect 61702 203630 61820 203690
rect 62806 203630 62908 203690
rect 63936 203690 63996 204000
rect 65296 203690 65356 204000
rect 66384 203690 66444 204000
rect 63936 203630 64154 203690
rect 51214 201245 51274 203630
rect 51211 201244 51277 201245
rect 51211 201180 51212 201244
rect 51276 201180 51277 201244
rect 51211 201179 51277 201180
rect 52318 200837 52378 203630
rect 53422 201245 53482 203630
rect 53419 201244 53485 201245
rect 53419 201180 53420 201244
rect 53484 201180 53485 201244
rect 53419 201179 53485 201180
rect 50107 200836 50173 200837
rect 50107 200772 50108 200836
rect 50172 200772 50173 200836
rect 50107 200771 50173 200772
rect 52315 200836 52381 200837
rect 52315 200772 52316 200836
rect 52380 200772 52381 200836
rect 52315 200771 52381 200772
rect 54526 200701 54586 203630
rect 55630 201245 55690 203630
rect 55794 201454 56414 202000
rect 55627 201244 55693 201245
rect 55627 201180 55628 201244
rect 55692 201180 55693 201244
rect 55627 201179 55693 201180
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 54523 200700 54589 200701
rect 54523 200636 54524 200700
rect 54588 200636 54589 200700
rect 54523 200635 54589 200636
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 165454 56414 200898
rect 56918 200701 56978 203630
rect 58022 201109 58082 203630
rect 59310 201245 59370 203630
rect 59307 201244 59373 201245
rect 59307 201180 59308 201244
rect 59372 201180 59373 201244
rect 59307 201179 59373 201180
rect 58019 201108 58085 201109
rect 58019 201044 58020 201108
rect 58084 201044 58085 201108
rect 58019 201043 58085 201044
rect 56915 200700 56981 200701
rect 56915 200636 56916 200700
rect 56980 200636 56981 200700
rect 56915 200635 56981 200636
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 169174 60134 202000
rect 60598 201109 60658 203630
rect 61702 201381 61762 203630
rect 61699 201380 61765 201381
rect 61699 201316 61700 201380
rect 61764 201316 61765 201380
rect 61699 201315 61765 201316
rect 62806 201245 62866 203630
rect 62803 201244 62869 201245
rect 62803 201180 62804 201244
rect 62868 201180 62869 201244
rect 62803 201179 62869 201180
rect 60595 201108 60661 201109
rect 60595 201044 60596 201108
rect 60660 201044 60661 201108
rect 60595 201043 60661 201044
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 172894 63854 202000
rect 64094 201381 64154 203630
rect 64646 203630 65356 203690
rect 66302 203630 66444 203690
rect 67608 203690 67668 204000
rect 68696 203690 68756 204000
rect 67608 203630 67834 203690
rect 64091 201380 64157 201381
rect 64091 201316 64092 201380
rect 64156 201316 64157 201380
rect 64091 201315 64157 201316
rect 64646 200293 64706 203630
rect 66302 200429 66362 203630
rect 66299 200428 66365 200429
rect 66299 200364 66300 200428
rect 66364 200364 66365 200428
rect 66299 200363 66365 200364
rect 64643 200292 64709 200293
rect 64643 200228 64644 200292
rect 64708 200228 64709 200292
rect 64643 200227 64709 200228
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 176614 67574 202000
rect 67774 200565 67834 203630
rect 68694 203630 68756 203690
rect 68694 201381 68754 203630
rect 69784 203557 69844 204000
rect 71144 203557 71204 204000
rect 72232 203557 72292 204000
rect 73320 203557 73380 204000
rect 74408 203557 74468 204000
rect 75768 203557 75828 204000
rect 76992 203690 77052 204000
rect 76974 203630 77052 203690
rect 69781 203556 69847 203557
rect 69781 203492 69782 203556
rect 69846 203492 69847 203556
rect 69781 203491 69847 203492
rect 71141 203556 71207 203557
rect 71141 203492 71142 203556
rect 71206 203492 71207 203556
rect 71141 203491 71207 203492
rect 72229 203556 72295 203557
rect 72229 203492 72230 203556
rect 72294 203492 72295 203556
rect 72229 203491 72295 203492
rect 73317 203556 73383 203557
rect 73317 203492 73318 203556
rect 73382 203492 73383 203556
rect 73317 203491 73383 203492
rect 74405 203556 74471 203557
rect 74405 203492 74406 203556
rect 74470 203492 74471 203556
rect 74405 203491 74471 203492
rect 75765 203556 75831 203557
rect 75765 203492 75766 203556
rect 75830 203492 75831 203556
rect 75765 203491 75831 203492
rect 76974 203013 77034 203630
rect 78080 203557 78140 204000
rect 79168 203690 79228 204000
rect 143224 203829 143284 204000
rect 143221 203828 143287 203829
rect 143221 203764 143222 203828
rect 143286 203764 143287 203828
rect 143221 203763 143287 203764
rect 143360 203690 143420 204000
rect 79168 203630 79242 203690
rect 143360 203630 143458 203690
rect 78077 203556 78143 203557
rect 78077 203492 78078 203556
rect 78142 203492 78143 203556
rect 78077 203491 78143 203492
rect 76971 203012 77037 203013
rect 76971 202948 76972 203012
rect 77036 202948 77037 203012
rect 76971 202947 77037 202948
rect 68691 201380 68757 201381
rect 68691 201316 68692 201380
rect 68756 201316 68757 201380
rect 68691 201315 68757 201316
rect 67771 200564 67837 200565
rect 67771 200500 67772 200564
rect 67836 200500 67837 200564
rect 67771 200499 67837 200500
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 183454 74414 202000
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 187174 78134 202000
rect 79182 201381 79242 203630
rect 79179 201380 79245 201381
rect 79179 201316 79180 201380
rect 79244 201316 79245 201380
rect 79179 201315 79245 201316
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 190894 81854 202000
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 194614 85574 202000
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 201454 92414 202000
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 169174 96134 202000
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 172894 99854 202000
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 176614 103574 202000
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 183454 110414 202000
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 187174 114134 202000
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 190894 117854 202000
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 194614 121574 202000
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 201454 128414 202000
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 169174 132134 202000
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 172894 135854 202000
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 176614 139574 202000
rect 143398 200837 143458 203630
rect 143395 200836 143461 200837
rect 143395 200772 143396 200836
rect 143460 200772 143461 200836
rect 143395 200771 143461 200772
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 183454 146414 202000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 187174 150134 202000
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 190894 153854 202000
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 194614 157574 202000
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 407708 182414 434898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 407708 186134 438618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 407708 189854 442338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 407708 193574 410058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 407708 200414 416898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 407708 204134 420618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 407708 207854 424338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 407708 211574 428058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 213499 408508 213565 408509
rect 213499 408444 213500 408508
rect 213564 408444 213565 408508
rect 213499 408443 213565 408444
rect 216259 408508 216325 408509
rect 216259 408444 216260 408508
rect 216324 408444 216325 408508
rect 216259 408443 216325 408444
rect 208715 407148 208781 407149
rect 208715 407084 208716 407148
rect 208780 407084 208781 407148
rect 208715 407083 208781 407084
rect 211107 407148 211173 407149
rect 211107 407084 211108 407148
rect 211172 407084 211173 407148
rect 211107 407083 211173 407084
rect 208718 406330 208778 407083
rect 211110 406330 211170 407083
rect 213502 406330 213562 408443
rect 216262 406330 216322 408443
rect 217794 407708 218414 434898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221043 408372 221109 408373
rect 221043 408308 221044 408372
rect 221108 408308 221109 408372
rect 221043 408307 221109 408308
rect 218467 407148 218533 407149
rect 218467 407084 218468 407148
rect 218532 407084 218533 407148
rect 218467 407083 218533 407084
rect 208704 406270 208778 406330
rect 211016 406270 211170 406330
rect 213464 406270 213562 406330
rect 216184 406270 216322 406330
rect 218470 406330 218530 407083
rect 221046 406330 221106 408307
rect 221514 407708 222134 438618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 223435 408372 223501 408373
rect 223435 408308 223436 408372
rect 223500 408308 223501 408372
rect 223435 408307 223501 408308
rect 223438 406330 223498 408307
rect 225234 407708 225854 442338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 239514 690600 240134 707162
rect 243234 690600 243854 709082
rect 246954 690600 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 690600 254414 704282
rect 257514 690600 258134 706202
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 690600 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 690600 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 690600 272414 705242
rect 275514 690600 276134 707162
rect 241080 687454 241480 687486
rect 241080 687218 241162 687454
rect 241398 687218 241480 687454
rect 241080 687134 241480 687218
rect 241080 686898 241162 687134
rect 241398 686898 241480 687134
rect 241080 686866 241480 686898
rect 243680 687454 244080 687486
rect 243680 687218 243762 687454
rect 243998 687218 244080 687454
rect 243680 687134 244080 687218
rect 243680 686898 243762 687134
rect 243998 686898 244080 687134
rect 243680 686866 244080 686898
rect 250880 687454 251280 687486
rect 250880 687218 250962 687454
rect 251198 687218 251280 687454
rect 250880 687134 251280 687218
rect 250880 686898 250962 687134
rect 251198 686898 251280 687134
rect 250880 686866 251280 686898
rect 258080 687454 258480 687486
rect 258080 687218 258162 687454
rect 258398 687218 258480 687454
rect 258080 687134 258480 687218
rect 258080 686898 258162 687134
rect 258398 686898 258480 687134
rect 258080 686866 258480 686898
rect 265280 687454 265680 687486
rect 265280 687218 265362 687454
rect 265598 687218 265680 687454
rect 265280 687134 265680 687218
rect 265280 686898 265362 687134
rect 265598 686898 265680 687134
rect 265280 686866 265680 686898
rect 272480 687454 272880 687486
rect 272480 687218 272562 687454
rect 272798 687218 272880 687454
rect 272480 687134 272880 687218
rect 272480 686898 272562 687134
rect 272798 686898 272880 687134
rect 272480 686866 272880 686898
rect 275080 687454 275480 687486
rect 275080 687218 275162 687454
rect 275398 687218 275480 687454
rect 275080 687134 275480 687218
rect 275080 686898 275162 687134
rect 275398 686898 275480 687134
rect 275080 686866 275480 686898
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 240080 669454 240480 669486
rect 240080 669218 240162 669454
rect 240398 669218 240480 669454
rect 240080 669134 240480 669218
rect 240080 668898 240162 669134
rect 240398 668898 240480 669134
rect 240080 668866 240480 668898
rect 247280 669454 247680 669486
rect 247280 669218 247362 669454
rect 247598 669218 247680 669454
rect 247280 669134 247680 669218
rect 247280 668898 247362 669134
rect 247598 668898 247680 669134
rect 247280 668866 247680 668898
rect 254480 669454 254880 669486
rect 254480 669218 254562 669454
rect 254798 669218 254880 669454
rect 254480 669134 254880 669218
rect 254480 668898 254562 669134
rect 254798 668898 254880 669134
rect 254480 668866 254880 668898
rect 261680 669454 262080 669486
rect 261680 669218 261762 669454
rect 261998 669218 262080 669454
rect 261680 669134 262080 669218
rect 261680 668898 261762 669134
rect 261998 668898 262080 669134
rect 261680 668866 262080 668898
rect 268880 669454 269280 669486
rect 268880 669218 268962 669454
rect 269198 669218 269280 669454
rect 268880 669134 269280 669218
rect 268880 668898 268962 669134
rect 269198 668898 269280 669134
rect 268880 668866 269280 668898
rect 276080 669454 276480 669486
rect 276080 669218 276162 669454
rect 276398 669218 276480 669454
rect 276080 669134 276480 669218
rect 276080 668898 276162 669134
rect 276398 668898 276480 669134
rect 276080 668866 276480 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 631820 236414 632898
rect 239514 637174 240134 665600
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 631820 240134 636618
rect 243234 640894 243854 665600
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 631820 243854 640338
rect 246954 644614 247574 665600
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 631820 247574 644058
rect 253794 651454 254414 665600
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 631820 254414 650898
rect 257514 655174 258134 665600
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 631820 258134 654618
rect 261234 658894 261854 665600
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 631820 261854 658338
rect 264954 662614 265574 665600
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 631820 265574 662058
rect 271794 633454 272414 665600
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 631820 272414 632898
rect 275514 637174 276134 665600
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 631820 276134 636618
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 631820 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 631820 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 631820 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 239408 615454 239728 615486
rect 239408 615218 239450 615454
rect 239686 615218 239728 615454
rect 239408 615134 239728 615218
rect 239408 614898 239450 615134
rect 239686 614898 239728 615134
rect 239408 614866 239728 614898
rect 270128 615454 270448 615486
rect 270128 615218 270170 615454
rect 270406 615218 270448 615454
rect 270128 615134 270448 615218
rect 270128 614898 270170 615134
rect 270406 614898 270448 615134
rect 270128 614866 270448 614898
rect 254768 597454 255088 597486
rect 254768 597218 254810 597454
rect 255046 597218 255088 597454
rect 254768 597134 255088 597218
rect 254768 596898 254810 597134
rect 255046 596898 255088 597134
rect 254768 596866 255088 596898
rect 285488 597454 285808 597486
rect 285488 597218 285530 597454
rect 285766 597218 285808 597454
rect 285488 597134 285808 597218
rect 285488 596898 285530 597134
rect 285766 596898 285808 597134
rect 285488 596866 285808 596898
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 239408 579454 239728 579486
rect 239408 579218 239450 579454
rect 239686 579218 239728 579454
rect 239408 579134 239728 579218
rect 239408 578898 239450 579134
rect 239686 578898 239728 579134
rect 239408 578866 239728 578898
rect 270128 579454 270448 579486
rect 270128 579218 270170 579454
rect 270406 579218 270448 579454
rect 270128 579134 270448 579218
rect 270128 578898 270170 579134
rect 270406 578898 270448 579134
rect 270128 578866 270448 578898
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 226195 408508 226261 408509
rect 226195 408444 226196 408508
rect 226260 408444 226261 408508
rect 226195 408443 226261 408444
rect 228587 408508 228653 408509
rect 228587 408444 228588 408508
rect 228652 408444 228653 408508
rect 228587 408443 228653 408444
rect 226198 406330 226258 408443
rect 228590 406330 228650 408443
rect 228954 407708 229574 410058
rect 235794 561454 236414 573820
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 407708 236414 416898
rect 239514 565174 240134 573820
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 407708 240134 420618
rect 243234 568894 243854 573820
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 407708 243854 424338
rect 246954 572614 247574 573820
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 407708 247574 428058
rect 253794 543454 254414 573820
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 251035 408508 251101 408509
rect 251035 408444 251036 408508
rect 251100 408444 251101 408508
rect 251035 408443 251101 408444
rect 253611 408508 253677 408509
rect 253611 408444 253612 408508
rect 253676 408444 253677 408508
rect 253611 408443 253677 408444
rect 231163 407148 231229 407149
rect 231163 407084 231164 407148
rect 231228 407084 231229 407148
rect 231163 407083 231229 407084
rect 233555 407148 233621 407149
rect 233555 407084 233556 407148
rect 233620 407084 233621 407148
rect 233555 407083 233621 407084
rect 236131 407148 236197 407149
rect 236131 407084 236132 407148
rect 236196 407084 236197 407148
rect 236131 407083 236197 407084
rect 240915 407148 240981 407149
rect 240915 407084 240916 407148
rect 240980 407084 240981 407148
rect 240915 407083 240981 407084
rect 246067 407148 246133 407149
rect 246067 407084 246068 407148
rect 246132 407084 246133 407148
rect 246067 407083 246133 407084
rect 248643 407148 248709 407149
rect 248643 407084 248644 407148
rect 248708 407084 248709 407148
rect 248643 407083 248709 407084
rect 231166 406330 231226 407083
rect 218470 406270 218556 406330
rect 221046 406270 221140 406330
rect 223438 406270 223588 406330
rect 208704 405620 208764 406270
rect 211016 405620 211076 406270
rect 213464 405620 213524 406270
rect 216184 405620 216244 406270
rect 218496 405620 218556 406270
rect 221080 405620 221140 406270
rect 223528 405620 223588 406270
rect 226112 406270 226258 406330
rect 228560 406270 228650 406330
rect 231144 406270 231226 406330
rect 233558 406330 233618 407083
rect 236134 406330 236194 407083
rect 238523 406604 238589 406605
rect 238523 406540 238524 406604
rect 238588 406540 238589 406604
rect 238523 406539 238589 406540
rect 238526 406330 238586 406539
rect 233558 406270 233652 406330
rect 236134 406270 236236 406330
rect 226112 405620 226172 406270
rect 228560 405620 228620 406270
rect 231144 405620 231204 406270
rect 233592 405620 233652 406270
rect 236176 405620 236236 406270
rect 238488 406270 238586 406330
rect 240918 406330 240978 407083
rect 243675 406604 243741 406605
rect 243675 406540 243676 406604
rect 243740 406540 243741 406604
rect 243675 406539 243741 406540
rect 243678 406330 243738 406539
rect 240918 406270 240996 406330
rect 238488 405620 238548 406270
rect 240936 405620 240996 406270
rect 243656 406270 243738 406330
rect 246070 406330 246130 407083
rect 248646 406330 248706 407083
rect 251038 406330 251098 408443
rect 253614 406330 253674 408443
rect 253794 407708 254414 434898
rect 257514 547174 258134 573820
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 407708 258134 438618
rect 261234 550894 261854 573820
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 258579 408508 258645 408509
rect 258579 408444 258580 408508
rect 258644 408444 258645 408508
rect 258579 408443 258645 408444
rect 256003 407148 256069 407149
rect 256003 407084 256004 407148
rect 256068 407084 256069 407148
rect 256003 407083 256069 407084
rect 256006 406330 256066 407083
rect 246070 406270 246164 406330
rect 243656 405620 243716 406270
rect 246104 405620 246164 406270
rect 248552 406270 248706 406330
rect 251000 406270 251098 406330
rect 253584 406270 253674 406330
rect 255896 406270 256066 406330
rect 258582 406330 258642 408443
rect 261234 407708 261854 442338
rect 264954 554614 265574 573820
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 263547 408508 263613 408509
rect 263547 408444 263548 408508
rect 263612 408444 263613 408508
rect 263547 408443 263613 408444
rect 261155 407148 261221 407149
rect 261155 407084 261156 407148
rect 261220 407084 261221 407148
rect 261155 407083 261221 407084
rect 261158 406330 261218 407083
rect 263550 406330 263610 408443
rect 264954 407708 265574 410058
rect 271794 561454 272414 573820
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 265939 408508 266005 408509
rect 265939 408444 265940 408508
rect 266004 408444 266005 408508
rect 265939 408443 266005 408444
rect 258582 406270 258676 406330
rect 248552 405620 248612 406270
rect 251000 405620 251060 406270
rect 253584 405620 253644 406270
rect 255896 405620 255956 406270
rect 258616 405620 258676 406270
rect 261064 406270 261218 406330
rect 263512 406270 263610 406330
rect 265942 406330 266002 408443
rect 271091 408372 271157 408373
rect 271091 408308 271092 408372
rect 271156 408308 271157 408372
rect 271091 408307 271157 408308
rect 268515 408100 268581 408101
rect 268515 408036 268516 408100
rect 268580 408036 268581 408100
rect 268515 408035 268581 408036
rect 268518 406330 268578 408035
rect 271094 406330 271154 408307
rect 271794 407708 272414 416898
rect 275514 565174 276134 573820
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 273667 408508 273733 408509
rect 273667 408444 273668 408508
rect 273732 408444 273733 408508
rect 273667 408443 273733 408444
rect 273670 406330 273730 408443
rect 275514 407708 276134 420618
rect 279234 568894 279854 573820
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 278451 408508 278517 408509
rect 278451 408444 278452 408508
rect 278516 408444 278517 408508
rect 278451 408443 278517 408444
rect 276059 407148 276125 407149
rect 276059 407084 276060 407148
rect 276124 407084 276125 407148
rect 276059 407083 276125 407084
rect 276062 406330 276122 407083
rect 265942 406270 266020 406330
rect 261064 405620 261124 406270
rect 263512 405620 263572 406270
rect 265960 405620 266020 406270
rect 268408 406270 268578 406330
rect 270992 406270 271154 406330
rect 273576 406270 273730 406330
rect 276024 406270 276122 406330
rect 278454 406330 278514 408443
rect 279234 407708 279854 424338
rect 282954 572614 283574 573820
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 407708 283574 428058
rect 289794 543454 290414 573820
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 286179 408372 286245 408373
rect 286179 408308 286180 408372
rect 286244 408308 286245 408372
rect 286179 408307 286245 408308
rect 283419 407148 283485 407149
rect 283419 407084 283420 407148
rect 283484 407084 283485 407148
rect 283419 407083 283485 407084
rect 281027 406604 281093 406605
rect 281027 406540 281028 406604
rect 281092 406540 281093 406604
rect 281027 406539 281093 406540
rect 281030 406330 281090 406539
rect 283422 406330 283482 407083
rect 286182 406330 286242 408307
rect 289794 407708 290414 434898
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 407708 294134 438618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 407708 297854 442338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 407708 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 407708 308414 416898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 407708 312134 420618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 407708 315854 424338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 298507 407148 298573 407149
rect 298507 407084 298508 407148
rect 298572 407084 298573 407148
rect 298507 407083 298573 407084
rect 299795 407148 299861 407149
rect 299795 407084 299796 407148
rect 299860 407084 299861 407148
rect 299795 407083 299861 407084
rect 310835 407148 310901 407149
rect 310835 407084 310836 407148
rect 310900 407084 310901 407148
rect 310835 407083 310901 407084
rect 298510 406330 298570 407083
rect 299798 406330 299858 407083
rect 278454 406270 278532 406330
rect 281030 406270 281116 406330
rect 268408 405620 268468 406270
rect 270992 405620 271052 406270
rect 273576 405620 273636 406270
rect 276024 405620 276084 406270
rect 278472 405620 278532 406270
rect 281056 405620 281116 406270
rect 283368 406270 283482 406330
rect 286088 406270 286242 406330
rect 298464 406270 298570 406330
rect 299688 406270 299858 406330
rect 310838 406330 310898 407083
rect 310838 406270 310900 406330
rect 283368 405620 283428 406270
rect 286088 405620 286148 406270
rect 298464 405620 298524 406270
rect 299688 405620 299748 406270
rect 310840 405620 310900 406270
rect 180952 399454 181300 399486
rect 180952 399218 181008 399454
rect 181244 399218 181300 399454
rect 180952 399134 181300 399218
rect 180952 398898 181008 399134
rect 181244 398898 181300 399134
rect 180952 398866 181300 398898
rect 315320 399454 315668 399486
rect 315320 399218 315376 399454
rect 315612 399218 315668 399454
rect 315320 399134 315668 399218
rect 315320 398898 315376 399134
rect 315612 398898 315668 399134
rect 315320 398866 315668 398898
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 180272 381454 180620 381486
rect 180272 381218 180328 381454
rect 180564 381218 180620 381454
rect 180272 381134 180620 381218
rect 180272 380898 180328 381134
rect 180564 380898 180620 381134
rect 180272 380866 180620 380898
rect 316000 381454 316348 381486
rect 316000 381218 316056 381454
rect 316292 381218 316348 381454
rect 316000 381134 316348 381218
rect 316000 380898 316056 381134
rect 316292 380898 316348 381134
rect 316000 380866 316348 380898
rect 180952 363454 181300 363486
rect 180952 363218 181008 363454
rect 181244 363218 181300 363454
rect 180952 363134 181300 363218
rect 180952 362898 181008 363134
rect 181244 362898 181300 363134
rect 180952 362866 181300 362898
rect 315320 363454 315668 363486
rect 315320 363218 315376 363454
rect 315612 363218 315668 363454
rect 315320 363134 315668 363218
rect 315320 362898 315376 363134
rect 315612 362898 315668 363134
rect 315320 362866 315668 362898
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 180272 345454 180620 345486
rect 180272 345218 180328 345454
rect 180564 345218 180620 345454
rect 180272 345134 180620 345218
rect 180272 344898 180328 345134
rect 180564 344898 180620 345134
rect 180272 344866 180620 344898
rect 316000 345454 316348 345486
rect 316000 345218 316056 345454
rect 316292 345218 316348 345454
rect 316000 345134 316348 345218
rect 316000 344898 316056 345134
rect 316292 344898 316348 345134
rect 316000 344866 316348 344898
rect 180952 327454 181300 327486
rect 180952 327218 181008 327454
rect 181244 327218 181300 327454
rect 180952 327134 181300 327218
rect 180952 326898 181008 327134
rect 181244 326898 181300 327134
rect 180952 326866 181300 326898
rect 315320 327454 315668 327486
rect 315320 327218 315376 327454
rect 315612 327218 315668 327454
rect 315320 327134 315668 327218
rect 315320 326898 315376 327134
rect 315612 326898 315668 327134
rect 315320 326866 315668 326898
rect 196056 322010 196116 322506
rect 197144 322010 197204 322506
rect 198232 322010 198292 322506
rect 199592 322010 199652 322506
rect 196022 321950 196116 322010
rect 197126 321950 197204 322010
rect 198230 321950 198292 322010
rect 199518 321950 199652 322010
rect 200544 322010 200604 322506
rect 201768 322010 201828 322506
rect 200544 321950 200682 322010
rect 179643 321876 179709 321877
rect 179643 321812 179644 321876
rect 179708 321812 179709 321876
rect 179643 321811 179709 321812
rect 179459 321740 179525 321741
rect 179459 321676 179460 321740
rect 179524 321676 179525 321740
rect 179459 321675 179525 321676
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 178539 320244 178605 320245
rect 178539 320180 178540 320244
rect 178604 320180 178605 320244
rect 178539 320179 178605 320180
rect 178723 320244 178789 320245
rect 178723 320180 178724 320244
rect 178788 320180 178789 320244
rect 178723 320179 178789 320180
rect 174954 301674 175574 320058
rect 177987 319156 178053 319157
rect 177987 319092 177988 319156
rect 178052 319092 178053 319156
rect 177987 319091 178053 319092
rect 177990 318885 178050 319091
rect 177987 318884 178053 318885
rect 177987 318820 177988 318884
rect 178052 318820 178053 318884
rect 177987 318819 178053 318820
rect 174954 301438 174986 301674
rect 175222 301438 175306 301674
rect 175542 301438 175574 301674
rect 174954 301354 175574 301438
rect 174954 301118 174986 301354
rect 175222 301118 175306 301354
rect 175542 301118 175574 301354
rect 174954 284614 175574 301118
rect 178355 288828 178421 288829
rect 178355 288764 178356 288828
rect 178420 288764 178421 288828
rect 178355 288763 178421 288764
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 178171 267748 178237 267749
rect 178171 267684 178172 267748
rect 178236 267684 178237 267748
rect 178171 267683 178237 267684
rect 178174 258229 178234 267683
rect 178171 258228 178237 258229
rect 178171 258164 178172 258228
rect 178236 258164 178237 258228
rect 178171 258163 178237 258164
rect 178171 257956 178237 257957
rect 178171 257892 178172 257956
rect 178236 257892 178237 257956
rect 178171 257891 178237 257892
rect 178174 253877 178234 257891
rect 178171 253876 178237 253877
rect 178171 253812 178172 253876
rect 178236 253812 178237 253876
rect 178171 253811 178237 253812
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 178358 244357 178418 288763
rect 178355 244356 178421 244357
rect 178355 244292 178356 244356
rect 178420 244292 178421 244356
rect 178355 244291 178421 244292
rect 178355 239460 178421 239461
rect 178355 239396 178356 239460
rect 178420 239396 178421 239460
rect 178355 239395 178421 239396
rect 178171 234428 178237 234429
rect 178171 234364 178172 234428
rect 178236 234364 178237 234428
rect 178171 234363 178237 234364
rect 178174 231870 178234 234363
rect 177990 231810 178234 231870
rect 177990 224773 178050 231810
rect 178171 224908 178237 224909
rect 178171 224844 178172 224908
rect 178236 224844 178237 224908
rect 178171 224843 178237 224844
rect 177987 224772 178053 224773
rect 177987 224708 177988 224772
rect 178052 224708 178053 224772
rect 177987 224707 178053 224708
rect 177803 222732 177869 222733
rect 177803 222668 177804 222732
rect 177868 222668 177869 222732
rect 177803 222667 177869 222668
rect 177806 215930 177866 222667
rect 178174 217290 178234 224843
rect 178358 220149 178418 239395
rect 178355 220148 178421 220149
rect 178355 220084 178356 220148
rect 178420 220084 178421 220148
rect 178355 220083 178421 220084
rect 178174 217230 178418 217290
rect 177806 215870 178234 215930
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 178174 205733 178234 215870
rect 178171 205732 178237 205733
rect 178171 205668 178172 205732
rect 178236 205668 178237 205732
rect 178171 205667 178237 205668
rect 178358 203149 178418 217230
rect 178355 203148 178421 203149
rect 178355 203084 178356 203148
rect 178420 203084 178421 203148
rect 178355 203083 178421 203084
rect 178542 201245 178602 320179
rect 178539 201244 178605 201245
rect 178539 201180 178540 201244
rect 178604 201180 178605 201244
rect 178539 201179 178605 201180
rect 178726 200293 178786 320179
rect 179275 319564 179341 319565
rect 179275 319500 179276 319564
rect 179340 319500 179341 319564
rect 179275 319499 179341 319500
rect 179091 319428 179157 319429
rect 179091 319364 179092 319428
rect 179156 319364 179157 319428
rect 179091 319363 179157 319364
rect 178907 319156 178973 319157
rect 178907 319092 178908 319156
rect 178972 319092 178973 319156
rect 178907 319091 178973 319092
rect 178910 200565 178970 319091
rect 178907 200564 178973 200565
rect 178907 200500 178908 200564
rect 178972 200500 178973 200564
rect 178907 200499 178973 200500
rect 178723 200292 178789 200293
rect 178723 200228 178724 200292
rect 178788 200228 178789 200292
rect 178723 200227 178789 200228
rect 179094 200157 179154 319363
rect 179278 288829 179338 319499
rect 179275 288828 179341 288829
rect 179275 288764 179276 288828
rect 179340 288764 179341 288828
rect 179275 288763 179341 288764
rect 179275 287876 179341 287877
rect 179275 287812 179276 287876
rect 179340 287812 179341 287876
rect 179275 287811 179341 287812
rect 179278 244629 179338 287811
rect 179275 244628 179341 244629
rect 179275 244564 179276 244628
rect 179340 244564 179341 244628
rect 179275 244563 179341 244564
rect 179275 244356 179341 244357
rect 179275 244292 179276 244356
rect 179340 244292 179341 244356
rect 179275 244291 179341 244292
rect 179278 239461 179338 244291
rect 179275 239460 179341 239461
rect 179275 239396 179276 239460
rect 179340 239396 179341 239460
rect 179275 239395 179341 239396
rect 179275 236604 179341 236605
rect 179275 236540 179276 236604
rect 179340 236540 179341 236604
rect 179275 236539 179341 236540
rect 179278 234837 179338 236539
rect 179275 234836 179341 234837
rect 179275 234772 179276 234836
rect 179340 234772 179341 234836
rect 179275 234771 179341 234772
rect 179275 234700 179341 234701
rect 179275 234636 179276 234700
rect 179340 234636 179341 234700
rect 179275 234635 179341 234636
rect 179278 234429 179338 234635
rect 179275 234428 179341 234429
rect 179275 234364 179276 234428
rect 179340 234364 179341 234428
rect 179275 234363 179341 234364
rect 179275 234292 179341 234293
rect 179275 234228 179276 234292
rect 179340 234228 179341 234292
rect 179275 234227 179341 234228
rect 179278 222733 179338 234227
rect 179462 233069 179522 321675
rect 179646 287877 179706 321811
rect 180011 321604 180077 321605
rect 180011 321540 180012 321604
rect 180076 321540 180077 321604
rect 180011 321539 180077 321540
rect 179827 320244 179893 320245
rect 179827 320180 179828 320244
rect 179892 320180 179893 320244
rect 179827 320179 179893 320180
rect 179643 287876 179709 287877
rect 179643 287812 179644 287876
rect 179708 287812 179709 287876
rect 179643 287811 179709 287812
rect 179643 287740 179709 287741
rect 179643 287676 179644 287740
rect 179708 287676 179709 287740
rect 179643 287675 179709 287676
rect 179646 244765 179706 287675
rect 179830 245989 179890 320179
rect 180014 287741 180074 321539
rect 180563 318884 180629 318885
rect 180563 318820 180564 318884
rect 180628 318820 180629 318884
rect 180563 318819 180629 318820
rect 180011 287740 180077 287741
rect 180011 287676 180012 287740
rect 180076 287676 180077 287740
rect 180011 287675 180077 287676
rect 180566 287469 180626 318819
rect 181794 291454 182414 320400
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 289308 182414 290898
rect 185514 295174 186134 320400
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 289308 186134 294618
rect 189234 298894 189854 320400
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 289308 189854 298338
rect 192954 302614 193574 320400
rect 196022 319429 196082 321950
rect 196019 319428 196085 319429
rect 196019 319364 196020 319428
rect 196084 319364 196085 319428
rect 196019 319363 196085 319364
rect 197126 318885 197186 321950
rect 198230 319429 198290 321950
rect 199518 319429 199578 321950
rect 198227 319428 198293 319429
rect 198227 319364 198228 319428
rect 198292 319364 198293 319428
rect 198227 319363 198293 319364
rect 199515 319428 199581 319429
rect 199515 319364 199516 319428
rect 199580 319364 199581 319428
rect 199515 319363 199581 319364
rect 197123 318884 197189 318885
rect 197123 318820 197124 318884
rect 197188 318820 197189 318884
rect 197123 318819 197189 318820
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 289308 193574 302058
rect 199794 309454 200414 320400
rect 200622 320109 200682 321950
rect 201726 321950 201828 322010
rect 203128 322010 203188 322506
rect 204216 322010 204276 322506
rect 205440 322010 205500 322506
rect 206528 322010 206588 322506
rect 207616 322010 207676 322506
rect 203128 321950 203258 322010
rect 204216 321950 204362 322010
rect 200619 320108 200685 320109
rect 200619 320044 200620 320108
rect 200684 320044 200685 320108
rect 200619 320043 200685 320044
rect 201726 319293 201786 321950
rect 203198 320109 203258 321950
rect 203195 320108 203261 320109
rect 203195 320044 203196 320108
rect 203260 320044 203261 320108
rect 203195 320043 203261 320044
rect 201723 319292 201789 319293
rect 201723 319228 201724 319292
rect 201788 319228 201789 319292
rect 201723 319227 201789 319228
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 289308 200414 308898
rect 203514 313174 204134 320400
rect 204302 320109 204362 321950
rect 205406 321950 205500 322010
rect 206510 321950 206588 322010
rect 207614 321950 207676 322010
rect 208704 322010 208764 322506
rect 210064 322010 210124 322506
rect 208704 321950 208778 322010
rect 204299 320108 204365 320109
rect 204299 320044 204300 320108
rect 204364 320044 204365 320108
rect 204299 320043 204365 320044
rect 205406 319157 205466 321950
rect 206510 319293 206570 321950
rect 207614 320653 207674 321950
rect 207611 320652 207677 320653
rect 207611 320588 207612 320652
rect 207676 320588 207677 320652
rect 207611 320587 207677 320588
rect 206507 319292 206573 319293
rect 206507 319228 206508 319292
rect 206572 319228 206573 319292
rect 206507 319227 206573 319228
rect 205403 319156 205469 319157
rect 205403 319092 205404 319156
rect 205468 319092 205469 319156
rect 205403 319091 205469 319092
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 289308 204134 312618
rect 207234 316894 207854 320400
rect 208718 319293 208778 321950
rect 210006 321950 210124 322010
rect 211288 322010 211348 322506
rect 212376 322010 212436 322506
rect 213464 322010 213524 322506
rect 214552 322010 214612 322506
rect 215912 322010 215972 322506
rect 217000 322010 217060 322506
rect 211288 321950 211722 322010
rect 212376 321950 212458 322010
rect 213464 321950 213562 322010
rect 214552 321950 214666 322010
rect 210006 319837 210066 321950
rect 210003 319836 210069 319837
rect 210003 319772 210004 319836
rect 210068 319772 210069 319836
rect 210003 319771 210069 319772
rect 208715 319292 208781 319293
rect 208715 319228 208716 319292
rect 208780 319228 208781 319292
rect 208715 319227 208781 319228
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 289308 207854 316338
rect 210954 301674 211574 320400
rect 211662 320109 211722 321950
rect 211659 320108 211725 320109
rect 211659 320044 211660 320108
rect 211724 320044 211725 320108
rect 211659 320043 211725 320044
rect 212398 319157 212458 321950
rect 213502 319429 213562 321950
rect 214606 319973 214666 321950
rect 215894 321950 215972 322010
rect 216998 321950 217060 322010
rect 218088 322010 218148 322506
rect 219448 322010 219508 322506
rect 218088 321950 218714 322010
rect 214603 319972 214669 319973
rect 214603 319908 214604 319972
rect 214668 319908 214669 319972
rect 214603 319907 214669 319908
rect 215894 319701 215954 321950
rect 216998 319701 217058 321950
rect 215891 319700 215957 319701
rect 215891 319636 215892 319700
rect 215956 319636 215957 319700
rect 215891 319635 215957 319636
rect 216995 319700 217061 319701
rect 216995 319636 216996 319700
rect 217060 319636 217061 319700
rect 216995 319635 217061 319636
rect 213499 319428 213565 319429
rect 213499 319364 213500 319428
rect 213564 319364 213565 319428
rect 213499 319363 213565 319364
rect 212395 319156 212461 319157
rect 212395 319092 212396 319156
rect 212460 319092 212461 319156
rect 212395 319091 212461 319092
rect 210954 301438 210986 301674
rect 211222 301438 211306 301674
rect 211542 301438 211574 301674
rect 210954 301354 211574 301438
rect 210954 301118 210986 301354
rect 211222 301118 211306 301354
rect 211542 301118 211574 301354
rect 208715 291140 208781 291141
rect 208715 291076 208716 291140
rect 208780 291076 208781 291140
rect 208715 291075 208781 291076
rect 210739 291140 210805 291141
rect 210739 291076 210740 291140
rect 210804 291076 210805 291140
rect 210739 291075 210805 291076
rect 208718 288010 208778 291075
rect 208704 287950 208778 288010
rect 210742 288010 210802 291075
rect 210954 289308 211574 301118
rect 217794 291454 218414 320400
rect 218654 319701 218714 321950
rect 219206 321950 219508 322010
rect 220672 322010 220732 322506
rect 221760 322010 221820 322506
rect 222848 322010 222908 322506
rect 223936 322010 223996 322506
rect 225296 322010 225356 322506
rect 226384 322010 226444 322506
rect 227608 322013 227668 322506
rect 228696 322013 228756 322506
rect 220672 321950 220738 322010
rect 221760 321950 221842 322010
rect 222848 321950 222946 322010
rect 223936 321950 224050 322010
rect 219206 321469 219266 321950
rect 220678 321469 220738 321950
rect 219203 321468 219269 321469
rect 219203 321404 219204 321468
rect 219268 321404 219269 321468
rect 219203 321403 219269 321404
rect 220675 321468 220741 321469
rect 220675 321404 220676 321468
rect 220740 321404 220741 321468
rect 220675 321403 220741 321404
rect 221782 320653 221842 321950
rect 221779 320652 221845 320653
rect 221779 320588 221780 320652
rect 221844 320588 221845 320652
rect 221779 320587 221845 320588
rect 218651 319700 218717 319701
rect 218651 319636 218652 319700
rect 218716 319636 218717 319700
rect 218651 319635 218717 319636
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 213499 291140 213565 291141
rect 213499 291076 213500 291140
rect 213564 291076 213565 291140
rect 213499 291075 213565 291076
rect 216259 291140 216325 291141
rect 216259 291076 216260 291140
rect 216324 291076 216325 291140
rect 216259 291075 216325 291076
rect 217794 291134 218414 291218
rect 221514 295174 222134 320400
rect 222886 319429 222946 321950
rect 223990 320109 224050 321950
rect 224910 321950 225356 322010
rect 226382 321950 226444 322010
rect 226931 322012 226997 322013
rect 223987 320108 224053 320109
rect 223987 320044 223988 320108
rect 224052 320044 224053 320108
rect 223987 320043 224053 320044
rect 222883 319428 222949 319429
rect 222883 319364 222884 319428
rect 222948 319364 222949 319428
rect 222883 319363 222949 319364
rect 224910 319293 224970 321950
rect 226382 321741 226442 321950
rect 226931 321948 226932 322012
rect 226996 321948 226997 322012
rect 226931 321947 226997 321948
rect 227605 322012 227671 322013
rect 227605 321948 227606 322012
rect 227670 321948 227671 322012
rect 227605 321947 227671 321948
rect 228693 322012 228759 322013
rect 228693 321948 228694 322012
rect 228758 321948 228759 322012
rect 229784 322010 229844 322506
rect 228693 321947 228759 321948
rect 229694 321950 229844 322010
rect 231144 322010 231204 322506
rect 232232 322010 232292 322506
rect 233350 322476 233434 322536
rect 231144 321950 231226 322010
rect 232232 321950 232330 322010
rect 226379 321740 226445 321741
rect 226379 321676 226380 321740
rect 226444 321676 226445 321740
rect 226379 321675 226445 321676
rect 224907 319292 224973 319293
rect 224907 319228 224908 319292
rect 224972 319228 224973 319292
rect 224907 319227 224973 319228
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 213502 288010 213562 291075
rect 216262 288010 216322 291075
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 218651 291140 218717 291141
rect 218651 291076 218652 291140
rect 218716 291076 218717 291140
rect 218651 291075 218717 291076
rect 221043 291140 221109 291141
rect 221043 291076 221044 291140
rect 221108 291076 221109 291140
rect 221043 291075 221109 291076
rect 217794 289308 218414 290898
rect 218654 288010 218714 291075
rect 210742 287950 211076 288010
rect 180563 287468 180629 287469
rect 180563 287404 180564 287468
rect 180628 287404 180629 287468
rect 180563 287403 180629 287404
rect 208704 287300 208764 287950
rect 211016 287300 211076 287950
rect 213464 287950 213562 288010
rect 216184 287950 216322 288010
rect 218496 287950 218714 288010
rect 221046 288010 221106 291075
rect 221514 289308 222134 294618
rect 225234 298894 225854 320400
rect 226382 320109 226442 321675
rect 226379 320108 226445 320109
rect 226379 320044 226380 320108
rect 226444 320044 226445 320108
rect 226379 320043 226445 320044
rect 226934 319973 226994 321947
rect 226931 319972 226997 319973
rect 226931 319908 226932 319972
rect 226996 319908 226997 319972
rect 226931 319907 226997 319908
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 223435 291140 223501 291141
rect 223435 291076 223436 291140
rect 223500 291076 223501 291140
rect 223435 291075 223501 291076
rect 223438 288010 223498 291075
rect 225234 289308 225854 298338
rect 228954 302614 229574 320400
rect 229694 319973 229754 321950
rect 231166 320109 231226 321950
rect 231163 320108 231229 320109
rect 231163 320044 231164 320108
rect 231228 320044 231229 320108
rect 231163 320043 231229 320044
rect 229691 319972 229757 319973
rect 229691 319908 229692 319972
rect 229756 319908 229757 319972
rect 229691 319907 229757 319908
rect 232270 319701 232330 321950
rect 232267 319700 232333 319701
rect 232267 319636 232268 319700
rect 232332 319636 232333 319700
rect 232267 319635 232333 319636
rect 233374 318885 233434 322476
rect 234408 322010 234468 322506
rect 235768 322010 235828 322506
rect 236992 322010 237052 322506
rect 238080 322010 238140 322506
rect 239168 322010 239228 322506
rect 303224 322010 303284 322506
rect 234294 321950 234468 322010
rect 235582 321950 235828 322010
rect 236870 321950 237052 322010
rect 237974 321950 238140 322010
rect 239078 321950 239228 322010
rect 303110 321950 303284 322010
rect 303360 322010 303420 322506
rect 303360 321950 303538 322010
rect 234294 319293 234354 321950
rect 235582 319293 235642 321950
rect 234291 319292 234357 319293
rect 234291 319228 234292 319292
rect 234356 319228 234357 319292
rect 234291 319227 234357 319228
rect 235579 319292 235645 319293
rect 235579 319228 235580 319292
rect 235644 319228 235645 319292
rect 235579 319227 235645 319228
rect 233371 318884 233437 318885
rect 233371 318820 233372 318884
rect 233436 318820 233437 318884
rect 233371 318819 233437 318820
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 226195 291140 226261 291141
rect 226195 291076 226196 291140
rect 226260 291076 226261 291140
rect 226195 291075 226261 291076
rect 228587 291140 228653 291141
rect 228587 291076 228588 291140
rect 228652 291076 228653 291140
rect 228587 291075 228653 291076
rect 226198 288010 226258 291075
rect 228590 288010 228650 291075
rect 228954 289308 229574 302058
rect 235794 309454 236414 320400
rect 236870 319565 236930 321950
rect 236867 319564 236933 319565
rect 236867 319500 236868 319564
rect 236932 319500 236933 319564
rect 236867 319499 236933 319500
rect 237974 319157 238034 321950
rect 237971 319156 238037 319157
rect 237971 319092 237972 319156
rect 238036 319092 238037 319156
rect 237971 319091 238037 319092
rect 239078 319021 239138 321950
rect 239075 319020 239141 319021
rect 239075 318956 239076 319020
rect 239140 318956 239141 319020
rect 239075 318955 239141 318956
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 231163 291140 231229 291141
rect 231163 291076 231164 291140
rect 231228 291076 231229 291140
rect 231163 291075 231229 291076
rect 231166 288010 231226 291075
rect 233555 290052 233621 290053
rect 233555 289988 233556 290052
rect 233620 289988 233621 290052
rect 233555 289987 233621 289988
rect 221046 287950 221140 288010
rect 223438 287950 223588 288010
rect 213464 287300 213524 287950
rect 216184 287300 216244 287950
rect 218496 287300 218556 287950
rect 221080 287300 221140 287950
rect 223528 287300 223588 287950
rect 226112 287950 226258 288010
rect 228560 287950 228650 288010
rect 231144 287950 231226 288010
rect 233558 288010 233618 289987
rect 235794 289308 236414 308898
rect 239514 313174 240134 320400
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 238523 291140 238589 291141
rect 238523 291076 238524 291140
rect 238588 291076 238589 291140
rect 238523 291075 238589 291076
rect 236499 291004 236565 291005
rect 236499 290940 236500 291004
rect 236564 290940 236565 291004
rect 236499 290939 236565 290940
rect 236502 288010 236562 290939
rect 238526 288010 238586 291075
rect 239514 289308 240134 312618
rect 243234 316894 243854 320400
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 240915 291140 240981 291141
rect 240915 291076 240916 291140
rect 240980 291076 240981 291140
rect 240915 291075 240981 291076
rect 233558 287950 233652 288010
rect 226112 287300 226172 287950
rect 228560 287300 228620 287950
rect 231144 287300 231204 287950
rect 233592 287300 233652 287950
rect 236176 287950 236562 288010
rect 238488 287950 238586 288010
rect 240918 288010 240978 291075
rect 243234 289308 243854 316338
rect 246954 301674 247574 320400
rect 246954 301438 246986 301674
rect 247222 301438 247306 301674
rect 247542 301438 247574 301674
rect 246954 301354 247574 301438
rect 246954 301118 246986 301354
rect 247222 301118 247306 301354
rect 247542 301118 247574 301354
rect 244043 291140 244109 291141
rect 244043 291076 244044 291140
rect 244108 291076 244109 291140
rect 244043 291075 244109 291076
rect 246067 291140 246133 291141
rect 246067 291076 246068 291140
rect 246132 291076 246133 291140
rect 246067 291075 246133 291076
rect 244046 288010 244106 291075
rect 240918 287950 240996 288010
rect 236176 287300 236236 287950
rect 238488 287300 238548 287950
rect 240936 287300 240996 287950
rect 243656 287950 244106 288010
rect 246070 288010 246130 291075
rect 246954 289308 247574 301118
rect 253794 291454 254414 320400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 248643 291140 248709 291141
rect 248643 291076 248644 291140
rect 248708 291076 248709 291140
rect 248643 291075 248709 291076
rect 251035 291140 251101 291141
rect 251035 291076 251036 291140
rect 251100 291076 251101 291140
rect 251035 291075 251101 291076
rect 253611 291140 253677 291141
rect 253611 291076 253612 291140
rect 253676 291076 253677 291140
rect 253611 291075 253677 291076
rect 253794 291134 254414 291218
rect 257514 295174 258134 320400
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 248646 288010 248706 291075
rect 251038 288010 251098 291075
rect 253614 288010 253674 291075
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 256003 291140 256069 291141
rect 256003 291076 256004 291140
rect 256068 291076 256069 291140
rect 256003 291075 256069 291076
rect 253794 289308 254414 290898
rect 256006 288010 256066 291075
rect 257514 289308 258134 294618
rect 261234 298894 261854 320400
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 258579 291140 258645 291141
rect 258579 291076 258580 291140
rect 258644 291076 258645 291140
rect 258579 291075 258645 291076
rect 246070 287950 246164 288010
rect 243656 287300 243716 287950
rect 246104 287300 246164 287950
rect 248552 287950 248706 288010
rect 251000 287950 251098 288010
rect 253584 287950 253674 288010
rect 255896 287950 256066 288010
rect 258582 288010 258642 291075
rect 260971 290460 261037 290461
rect 260971 290396 260972 290460
rect 261036 290396 261037 290460
rect 260971 290395 261037 290396
rect 260974 288010 261034 290395
rect 261234 289308 261854 298338
rect 264954 302614 265574 320400
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 263547 291140 263613 291141
rect 263547 291076 263548 291140
rect 263612 291076 263613 291140
rect 263547 291075 263613 291076
rect 263550 288010 263610 291075
rect 264954 289308 265574 302058
rect 271794 309454 272414 320400
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 268515 291140 268581 291141
rect 268515 291076 268516 291140
rect 268580 291076 268581 291140
rect 268515 291075 268581 291076
rect 271091 291140 271157 291141
rect 271091 291076 271092 291140
rect 271156 291076 271157 291140
rect 271091 291075 271157 291076
rect 265939 290732 266005 290733
rect 265939 290668 265940 290732
rect 266004 290668 266005 290732
rect 265939 290667 266005 290668
rect 258582 287950 258676 288010
rect 260974 287950 261124 288010
rect 248552 287300 248612 287950
rect 251000 287300 251060 287950
rect 253584 287300 253644 287950
rect 255896 287300 255956 287950
rect 258616 287300 258676 287950
rect 261064 287300 261124 287950
rect 263512 287950 263610 288010
rect 265942 288010 266002 290667
rect 268518 288010 268578 291075
rect 271094 288010 271154 291075
rect 271794 289308 272414 308898
rect 275514 313174 276134 320400
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 273667 291140 273733 291141
rect 273667 291076 273668 291140
rect 273732 291076 273733 291140
rect 273667 291075 273733 291076
rect 273670 288010 273730 291075
rect 275514 289308 276134 312618
rect 279234 316894 279854 320400
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 276243 291140 276309 291141
rect 276243 291076 276244 291140
rect 276308 291076 276309 291140
rect 276243 291075 276309 291076
rect 276246 288010 276306 291075
rect 277347 290732 277413 290733
rect 277347 290730 277348 290732
rect 265942 287950 266020 288010
rect 263512 287300 263572 287950
rect 265960 287300 266020 287950
rect 268408 287950 268578 288010
rect 270992 287950 271154 288010
rect 273576 287950 273730 288010
rect 276024 287950 276306 288010
rect 277166 290670 277348 290730
rect 277166 288010 277226 290670
rect 277347 290668 277348 290670
rect 277412 290668 277413 290732
rect 277347 290667 277413 290668
rect 279234 289308 279854 316338
rect 282954 301674 283574 320400
rect 282954 301438 282986 301674
rect 283222 301438 283306 301674
rect 283542 301438 283574 301674
rect 282954 301354 283574 301438
rect 282954 301118 282986 301354
rect 283222 301118 283306 301354
rect 283542 301118 283574 301354
rect 281027 291140 281093 291141
rect 281027 291076 281028 291140
rect 281092 291076 281093 291140
rect 281027 291075 281093 291076
rect 281030 288010 281090 291075
rect 282954 289308 283574 301118
rect 289794 291454 290414 320400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 283787 291140 283853 291141
rect 283787 291076 283788 291140
rect 283852 291076 283853 291140
rect 283787 291075 283853 291076
rect 289794 291134 290414 291218
rect 283790 288010 283850 291075
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 286179 289916 286245 289917
rect 286179 289852 286180 289916
rect 286244 289852 286245 289916
rect 286179 289851 286245 289852
rect 286182 288010 286242 289851
rect 289794 289308 290414 290898
rect 293514 295174 294134 320400
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 289308 294134 294618
rect 297234 298894 297854 320400
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 289308 297854 298338
rect 300954 302614 301574 320400
rect 303110 319429 303170 321950
rect 303107 319428 303173 319429
rect 303107 319364 303108 319428
rect 303172 319364 303173 319428
rect 303107 319363 303173 319364
rect 303478 319293 303538 321950
rect 318954 320614 319574 356058
rect 303475 319292 303541 319293
rect 303475 319228 303476 319292
rect 303540 319228 303541 319292
rect 303475 319227 303541 319228
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 298507 289916 298573 289917
rect 298507 289852 298508 289916
rect 298572 289852 298573 289916
rect 298507 289851 298573 289852
rect 299611 289916 299677 289917
rect 299611 289852 299612 289916
rect 299676 289852 299677 289916
rect 299611 289851 299677 289852
rect 298510 288010 298570 289851
rect 277166 287950 278532 288010
rect 281030 287950 281116 288010
rect 268408 287300 268468 287950
rect 270992 287300 271052 287950
rect 273576 287300 273636 287950
rect 276024 287300 276084 287950
rect 278472 287300 278532 287950
rect 281056 287300 281116 287950
rect 283368 287950 283850 288010
rect 286088 287950 286242 288010
rect 298464 287950 298570 288010
rect 299614 288010 299674 289851
rect 300954 289308 301574 302058
rect 307794 309454 308414 320400
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 289308 308414 308898
rect 311514 313174 312134 320400
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 310835 289916 310901 289917
rect 310835 289852 310836 289916
rect 310900 289852 310901 289916
rect 310835 289851 310901 289852
rect 310838 288010 310898 289851
rect 311514 289308 312134 312618
rect 315234 316894 315854 320400
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 289308 315854 316338
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 299614 287950 299748 288010
rect 310838 287950 310900 288010
rect 283368 287300 283428 287950
rect 286088 287300 286148 287950
rect 298464 287300 298524 287950
rect 299688 287300 299748 287950
rect 310840 287300 310900 287950
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 180272 273454 180620 273486
rect 180272 273218 180328 273454
rect 180564 273218 180620 273454
rect 180272 273134 180620 273218
rect 180272 272898 180328 273134
rect 180564 272898 180620 273134
rect 180272 272866 180620 272898
rect 316000 273454 316348 273486
rect 316000 273218 316056 273454
rect 316292 273218 316348 273454
rect 316000 273134 316348 273218
rect 316000 272898 316056 273134
rect 316292 272898 316348 273134
rect 316000 272866 316348 272898
rect 180952 255454 181300 255486
rect 180952 255218 181008 255454
rect 181244 255218 181300 255454
rect 180952 255134 181300 255218
rect 180952 254898 181008 255134
rect 181244 254898 181300 255134
rect 180952 254866 181300 254898
rect 315320 255454 315668 255486
rect 315320 255218 315376 255454
rect 315612 255218 315668 255454
rect 315320 255134 315668 255218
rect 315320 254898 315376 255134
rect 315612 254898 315668 255134
rect 315320 254866 315668 254898
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 179827 245988 179893 245989
rect 179827 245924 179828 245988
rect 179892 245924 179893 245988
rect 179827 245923 179893 245924
rect 179827 245716 179893 245717
rect 179827 245652 179828 245716
rect 179892 245652 179893 245716
rect 179827 245651 179893 245652
rect 179643 244764 179709 244765
rect 179643 244700 179644 244764
rect 179708 244700 179709 244764
rect 179643 244699 179709 244700
rect 179643 244356 179709 244357
rect 179643 244292 179644 244356
rect 179708 244292 179709 244356
rect 179643 244291 179709 244292
rect 179646 243949 179706 244291
rect 179830 243949 179890 245651
rect 179643 243948 179709 243949
rect 179643 243884 179644 243948
rect 179708 243884 179709 243948
rect 179643 243883 179709 243884
rect 179827 243948 179893 243949
rect 179827 243884 179828 243948
rect 179892 243884 179893 243948
rect 179827 243883 179893 243884
rect 179643 243812 179709 243813
rect 179643 243748 179644 243812
rect 179708 243748 179709 243812
rect 179643 243747 179709 243748
rect 179646 236605 179706 243747
rect 179827 243676 179893 243677
rect 179827 243612 179828 243676
rect 179892 243612 179893 243676
rect 179827 243611 179893 243612
rect 179643 236604 179709 236605
rect 179643 236540 179644 236604
rect 179708 236540 179709 236604
rect 179643 236539 179709 236540
rect 179643 236468 179709 236469
rect 179643 236404 179644 236468
rect 179708 236404 179709 236468
rect 179643 236403 179709 236404
rect 179646 233069 179706 236403
rect 179830 235650 179890 243611
rect 180272 237454 180620 237486
rect 180272 237218 180328 237454
rect 180564 237218 180620 237454
rect 180272 237134 180620 237218
rect 180272 236898 180328 237134
rect 180564 236898 180620 237134
rect 180272 236866 180620 236898
rect 316000 237454 316348 237486
rect 316000 237218 316056 237454
rect 316292 237218 316348 237454
rect 316000 237134 316348 237218
rect 316000 236898 316056 237134
rect 316292 236898 316348 237134
rect 316000 236866 316348 236898
rect 179830 235590 180062 235650
rect 180002 234834 180062 235590
rect 179830 234774 180062 234834
rect 179830 233069 179890 234774
rect 179459 233068 179525 233069
rect 179459 233004 179460 233068
rect 179524 233004 179525 233068
rect 179459 233003 179525 233004
rect 179643 233068 179709 233069
rect 179643 233004 179644 233068
rect 179708 233004 179709 233068
rect 179643 233003 179709 233004
rect 179827 233068 179893 233069
rect 179827 233004 179828 233068
rect 179892 233004 179893 233068
rect 179827 233003 179893 233004
rect 179459 232796 179525 232797
rect 179459 232732 179460 232796
rect 179524 232732 179525 232796
rect 179459 232731 179525 232732
rect 179643 232796 179709 232797
rect 179643 232732 179644 232796
rect 179708 232732 179709 232796
rect 179643 232731 179709 232732
rect 179827 232796 179893 232797
rect 179827 232732 179828 232796
rect 179892 232732 179893 232796
rect 179827 232731 179893 232732
rect 179462 224909 179522 232731
rect 179646 224909 179706 232731
rect 179830 225450 179890 232731
rect 179830 225390 180062 225450
rect 179459 224908 179525 224909
rect 179459 224844 179460 224908
rect 179524 224844 179525 224908
rect 179459 224843 179525 224844
rect 179643 224908 179709 224909
rect 179643 224844 179644 224908
rect 179708 224844 179709 224908
rect 179643 224843 179709 224844
rect 179459 224772 179525 224773
rect 179459 224708 179460 224772
rect 179524 224708 179525 224772
rect 179459 224707 179525 224708
rect 179275 222732 179341 222733
rect 179275 222668 179276 222732
rect 179340 222668 179341 222732
rect 179275 222667 179341 222668
rect 179275 220148 179341 220149
rect 179275 220084 179276 220148
rect 179340 220084 179341 220148
rect 179275 220083 179341 220084
rect 179278 200837 179338 220083
rect 179462 205869 179522 224707
rect 179643 224636 179709 224637
rect 179643 224572 179644 224636
rect 179708 224572 179709 224636
rect 180002 224634 180062 225390
rect 179643 224571 179709 224572
rect 179830 224574 180062 224634
rect 179646 210490 179706 224571
rect 179830 210629 179890 224574
rect 180952 219454 181300 219486
rect 180952 219218 181008 219454
rect 181244 219218 181300 219454
rect 180952 219134 181300 219218
rect 180952 218898 181008 219134
rect 181244 218898 181300 219134
rect 180952 218866 181300 218898
rect 315320 219454 315668 219486
rect 315320 219218 315376 219454
rect 315612 219218 315668 219454
rect 315320 219134 315668 219218
rect 315320 218898 315376 219134
rect 315612 218898 315668 219134
rect 315320 218866 315668 218898
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 179827 210628 179893 210629
rect 179827 210564 179828 210628
rect 179892 210564 179893 210628
rect 179827 210563 179893 210564
rect 179646 210430 179890 210490
rect 179643 210356 179709 210357
rect 179643 210292 179644 210356
rect 179708 210292 179709 210356
rect 179643 210291 179709 210292
rect 179459 205868 179525 205869
rect 179459 205804 179460 205868
rect 179524 205804 179525 205868
rect 179459 205803 179525 205804
rect 179646 205730 179706 210291
rect 179462 205670 179706 205730
rect 179462 201109 179522 205670
rect 179643 205596 179709 205597
rect 179643 205532 179644 205596
rect 179708 205532 179709 205596
rect 179643 205531 179709 205532
rect 179646 203285 179706 205531
rect 179643 203284 179709 203285
rect 179643 203220 179644 203284
rect 179708 203220 179709 203284
rect 179643 203219 179709 203220
rect 179830 203013 179890 210430
rect 180011 203828 180077 203829
rect 180011 203764 180012 203828
rect 180076 203764 180077 203828
rect 180011 203763 180077 203764
rect 179827 203012 179893 203013
rect 179827 202948 179828 203012
rect 179892 202948 179893 203012
rect 179827 202947 179893 202948
rect 179459 201108 179525 201109
rect 179459 201044 179460 201108
rect 179524 201044 179525 201108
rect 179459 201043 179525 201044
rect 180014 200973 180074 203763
rect 196056 203690 196116 204000
rect 197144 203690 197204 204000
rect 198232 203690 198292 204000
rect 199592 203690 199652 204000
rect 196022 203630 196116 203690
rect 197126 203630 197204 203690
rect 198230 203630 198292 203690
rect 199518 203630 199652 203690
rect 180011 200972 180077 200973
rect 180011 200908 180012 200972
rect 180076 200908 180077 200972
rect 180011 200907 180077 200908
rect 179275 200836 179341 200837
rect 179275 200772 179276 200836
rect 179340 200772 179341 200836
rect 179275 200771 179341 200772
rect 179091 200156 179157 200157
rect 179091 200092 179092 200156
rect 179156 200092 179157 200156
rect 179091 200091 179157 200092
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 183454 182414 202000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 187174 186134 202000
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 190894 189854 202000
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 194614 193574 202000
rect 196022 201381 196082 203630
rect 197126 201381 197186 203630
rect 198230 201381 198290 203630
rect 199518 201381 199578 203630
rect 200544 203554 200604 204000
rect 201768 203554 201828 204000
rect 203128 203554 203188 204000
rect 200544 203494 200682 203554
rect 199794 201454 200414 202000
rect 196019 201380 196085 201381
rect 196019 201316 196020 201380
rect 196084 201316 196085 201380
rect 196019 201315 196085 201316
rect 197123 201380 197189 201381
rect 197123 201316 197124 201380
rect 197188 201316 197189 201380
rect 197123 201315 197189 201316
rect 198227 201380 198293 201381
rect 198227 201316 198228 201380
rect 198292 201316 198293 201380
rect 198227 201315 198293 201316
rect 199515 201380 199581 201381
rect 199515 201316 199516 201380
rect 199580 201316 199581 201380
rect 199515 201315 199581 201316
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 200622 201381 200682 203494
rect 201726 203494 201828 203554
rect 203014 203494 203188 203554
rect 204216 203554 204276 204000
rect 205440 203554 205500 204000
rect 206528 203554 206588 204000
rect 207616 203554 207676 204000
rect 204216 203494 204362 203554
rect 200619 201380 200685 201381
rect 200619 201316 200620 201380
rect 200684 201316 200685 201380
rect 200619 201315 200685 201316
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 201726 200565 201786 203494
rect 203014 201245 203074 203494
rect 203011 201244 203077 201245
rect 203011 201180 203012 201244
rect 203076 201180 203077 201244
rect 203011 201179 203077 201180
rect 201723 200564 201789 200565
rect 201723 200500 201724 200564
rect 201788 200500 201789 200564
rect 201723 200499 201789 200500
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 202000
rect 204302 201245 204362 203494
rect 205406 203494 205500 203554
rect 206510 203494 206588 203554
rect 207062 203494 207676 203554
rect 208704 203554 208764 204000
rect 210064 203554 210124 204000
rect 208704 203494 208778 203554
rect 205406 201381 205466 203494
rect 205403 201380 205469 201381
rect 205403 201316 205404 201380
rect 205468 201316 205469 201380
rect 205403 201315 205469 201316
rect 204299 201244 204365 201245
rect 204299 201180 204300 201244
rect 204364 201180 204365 201244
rect 204299 201179 204365 201180
rect 206510 200157 206570 203494
rect 207062 200565 207122 203494
rect 207059 200564 207125 200565
rect 207059 200500 207060 200564
rect 207124 200500 207125 200564
rect 207059 200499 207125 200500
rect 206507 200156 206573 200157
rect 206507 200092 206508 200156
rect 206572 200092 206573 200156
rect 206507 200091 206573 200092
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 172894 207854 202000
rect 208718 200837 208778 203494
rect 210006 203494 210124 203554
rect 211288 203554 211348 204000
rect 212376 203554 212436 204000
rect 213464 203554 213524 204000
rect 214552 203554 214612 204000
rect 215912 203554 215972 204000
rect 217000 203554 217060 204000
rect 211288 203494 211722 203554
rect 212376 203494 212458 203554
rect 213464 203494 213562 203554
rect 214552 203494 214666 203554
rect 210006 200837 210066 203494
rect 208715 200836 208781 200837
rect 208715 200772 208716 200836
rect 208780 200772 208781 200836
rect 208715 200771 208781 200772
rect 210003 200836 210069 200837
rect 210003 200772 210004 200836
rect 210068 200772 210069 200836
rect 210003 200771 210069 200772
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 202000
rect 211662 201381 211722 203494
rect 211659 201380 211725 201381
rect 211659 201316 211660 201380
rect 211724 201316 211725 201380
rect 211659 201315 211725 201316
rect 212398 201109 212458 203494
rect 212395 201108 212461 201109
rect 212395 201044 212396 201108
rect 212460 201044 212461 201108
rect 212395 201043 212461 201044
rect 213502 200973 213562 203494
rect 214606 201245 214666 203494
rect 215894 203494 215972 203554
rect 216998 203494 217060 203554
rect 218088 203554 218148 204000
rect 219448 203690 219508 204000
rect 220672 203690 220732 204000
rect 221760 203690 221820 204000
rect 219448 203630 219634 203690
rect 220672 203630 220738 203690
rect 218088 203494 218714 203554
rect 215894 201245 215954 203494
rect 214603 201244 214669 201245
rect 214603 201180 214604 201244
rect 214668 201180 214669 201244
rect 214603 201179 214669 201180
rect 215891 201244 215957 201245
rect 215891 201180 215892 201244
rect 215956 201180 215957 201244
rect 215891 201179 215957 201180
rect 213499 200972 213565 200973
rect 213499 200908 213500 200972
rect 213564 200908 213565 200972
rect 213499 200907 213565 200908
rect 216998 200293 217058 203494
rect 216995 200292 217061 200293
rect 216995 200228 216996 200292
rect 217060 200228 217061 200292
rect 216995 200227 217061 200228
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 183454 218414 202000
rect 218654 200429 218714 203494
rect 219574 201245 219634 203630
rect 220678 201381 220738 203630
rect 221230 203630 221820 203690
rect 222848 203690 222908 204000
rect 223936 203690 223996 204000
rect 225296 203690 225356 204000
rect 226384 203690 226444 204000
rect 227608 203690 227668 204000
rect 228696 203690 228756 204000
rect 222848 203630 222946 203690
rect 223936 203630 224050 203690
rect 220675 201380 220741 201381
rect 220675 201316 220676 201380
rect 220740 201316 220741 201380
rect 220675 201315 220741 201316
rect 219571 201244 219637 201245
rect 219571 201180 219572 201244
rect 219636 201180 219637 201244
rect 219571 201179 219637 201180
rect 218651 200428 218717 200429
rect 218651 200364 218652 200428
rect 218716 200364 218717 200428
rect 218651 200363 218717 200364
rect 221230 200293 221290 203630
rect 221227 200292 221293 200293
rect 221227 200228 221228 200292
rect 221292 200228 221293 200292
rect 221227 200227 221293 200228
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 187174 222134 202000
rect 222886 201381 222946 203630
rect 223990 201381 224050 203630
rect 224910 203630 225356 203690
rect 226382 203630 226444 203690
rect 227486 203630 227668 203690
rect 228590 203630 228756 203690
rect 224910 201381 224970 203630
rect 226382 203149 226442 203630
rect 227486 203285 227546 203630
rect 227483 203284 227549 203285
rect 227483 203220 227484 203284
rect 227548 203220 227549 203284
rect 227483 203219 227549 203220
rect 226379 203148 226445 203149
rect 226379 203084 226380 203148
rect 226444 203084 226445 203148
rect 226379 203083 226445 203084
rect 228590 203013 228650 203630
rect 229784 203557 229844 204000
rect 231144 203557 231204 204000
rect 232232 203557 232292 204000
rect 233320 203557 233380 204000
rect 234408 203557 234468 204000
rect 235768 203557 235828 204000
rect 236992 203557 237052 204000
rect 238080 203557 238140 204000
rect 239168 203690 239228 204000
rect 303224 203690 303284 204000
rect 238526 203630 239228 203690
rect 303110 203630 303284 203690
rect 303360 203690 303420 204000
rect 303360 203630 303538 203690
rect 229781 203556 229847 203557
rect 229781 203492 229782 203556
rect 229846 203492 229847 203556
rect 229781 203491 229847 203492
rect 231141 203556 231207 203557
rect 231141 203492 231142 203556
rect 231206 203492 231207 203556
rect 231141 203491 231207 203492
rect 232229 203556 232295 203557
rect 232229 203492 232230 203556
rect 232294 203492 232295 203556
rect 232229 203491 232295 203492
rect 233317 203556 233383 203557
rect 233317 203492 233318 203556
rect 233382 203492 233383 203556
rect 233317 203491 233383 203492
rect 234405 203556 234471 203557
rect 234405 203492 234406 203556
rect 234470 203492 234471 203556
rect 234405 203491 234471 203492
rect 235765 203556 235831 203557
rect 235765 203492 235766 203556
rect 235830 203492 235831 203556
rect 235765 203491 235831 203492
rect 236989 203556 237055 203557
rect 236989 203492 236990 203556
rect 237054 203492 237055 203556
rect 236989 203491 237055 203492
rect 238077 203556 238143 203557
rect 238077 203492 238078 203556
rect 238142 203492 238143 203556
rect 238077 203491 238143 203492
rect 228587 203012 228653 203013
rect 228587 202948 228588 203012
rect 228652 202948 228653 203012
rect 228587 202947 228653 202948
rect 222883 201380 222949 201381
rect 222883 201316 222884 201380
rect 222948 201316 222949 201380
rect 222883 201315 222949 201316
rect 223987 201380 224053 201381
rect 223987 201316 223988 201380
rect 224052 201316 224053 201380
rect 223987 201315 224053 201316
rect 224907 201380 224973 201381
rect 224907 201316 224908 201380
rect 224972 201316 224973 201380
rect 224907 201315 224973 201316
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 190894 225854 202000
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 194614 229574 202000
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 201454 236414 202000
rect 238526 201650 238586 203630
rect 238526 201590 238954 201650
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 238894 201381 238954 201590
rect 238891 201380 238957 201381
rect 238891 201316 238892 201380
rect 238956 201316 238957 201380
rect 238891 201315 238957 201316
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 169174 240134 202000
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 202000
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 202000
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 183454 254414 202000
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 202000
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 202000
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 202000
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 201454 272414 202000
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 202000
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 202000
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 176614 283574 202000
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 183454 290414 202000
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 187174 294134 202000
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 190894 297854 202000
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 194614 301574 202000
rect 303110 201381 303170 203630
rect 303478 201381 303538 203630
rect 307794 201454 308414 202000
rect 303107 201380 303173 201381
rect 303107 201316 303108 201380
rect 303172 201316 303173 201380
rect 303107 201315 303173 201316
rect 303475 201380 303541 201381
rect 303475 201316 303476 201380
rect 303540 201316 303541 201380
rect 303475 201315 303541 201316
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 202000
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 202000
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 400000 344414 416898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 400000 348134 420618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 400000 351854 424338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 400000 355574 428058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 400000 362414 434898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 400000 366134 402618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 400000 369854 406338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 400000 373574 410058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 400000 380414 416898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 400000 384134 420618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 400000 387854 424338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 400000 391574 428058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 400000 398414 434898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 400000 402134 402618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 400000 405854 406338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 400000 409574 410058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 400000 416414 416898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 400000 420134 420618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 400000 423854 424338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 400000 427574 428058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 400000 434414 434898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 400000 438134 402618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 400000 441854 406338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 400000 445574 410058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 400000 452414 416898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 400000 456134 420618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 400000 459854 424338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 400000 463574 428058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 631820 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 631820 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 690600 488414 705242
rect 491514 690600 492134 707162
rect 495234 690600 495854 709082
rect 498954 690600 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 690600 506414 704282
rect 509514 690600 510134 706202
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 486240 687454 486640 687486
rect 486240 687218 486322 687454
rect 486558 687218 486640 687454
rect 486240 687134 486640 687218
rect 486240 686898 486322 687134
rect 486558 686898 486640 687134
rect 486240 686866 486640 686898
rect 489840 687454 490240 687486
rect 489840 687218 489922 687454
rect 490158 687218 490240 687454
rect 489840 687134 490240 687218
rect 489840 686898 489922 687134
rect 490158 686898 490240 687134
rect 489840 686866 490240 686898
rect 495440 687454 495840 687486
rect 495440 687218 495522 687454
rect 495758 687218 495840 687454
rect 495440 687134 495840 687218
rect 495440 686898 495522 687134
rect 495758 686898 495840 687134
rect 495440 686866 495840 686898
rect 501040 687454 501440 687486
rect 501040 687218 501122 687454
rect 501358 687218 501440 687454
rect 501040 687134 501440 687218
rect 501040 686898 501122 687134
rect 501358 686898 501440 687134
rect 501040 686866 501440 686898
rect 506640 687454 507040 687486
rect 506640 687218 506722 687454
rect 506958 687218 507040 687454
rect 506640 687134 507040 687218
rect 506640 686898 506722 687134
rect 506958 686898 507040 687134
rect 506640 686866 507040 686898
rect 510240 687454 510640 687486
rect 510240 687218 510322 687454
rect 510558 687218 510640 687454
rect 510240 687134 510640 687218
rect 510240 686898 510322 687134
rect 510558 686898 510640 687134
rect 510240 686866 510640 686898
rect 487040 669454 487440 669486
rect 487040 669218 487122 669454
rect 487358 669218 487440 669454
rect 487040 669134 487440 669218
rect 487040 668898 487122 669134
rect 487358 668898 487440 669134
rect 487040 668866 487440 668898
rect 492640 669454 493040 669486
rect 492640 669218 492722 669454
rect 492958 669218 493040 669454
rect 492640 669134 493040 669218
rect 492640 668898 492722 669134
rect 492958 668898 493040 669134
rect 492640 668866 493040 668898
rect 498240 669454 498640 669486
rect 498240 669218 498322 669454
rect 498558 669218 498640 669454
rect 498240 669134 498640 669218
rect 498240 668898 498322 669134
rect 498558 668898 498640 669134
rect 498240 668866 498640 668898
rect 503840 669454 504240 669486
rect 503840 669218 503922 669454
rect 504158 669218 504240 669454
rect 503840 669134 504240 669218
rect 503840 668898 503922 669134
rect 504158 668898 504240 669134
rect 503840 668866 504240 668898
rect 509440 669454 509840 669486
rect 509440 669218 509522 669454
rect 509758 669218 509840 669454
rect 509440 669134 509840 669218
rect 509440 668898 509522 669134
rect 509758 668898 509840 669134
rect 509440 668866 509840 668898
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 631820 481574 662058
rect 487794 633454 488414 665600
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 631820 488414 632898
rect 491514 637174 492134 665600
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 631820 492134 636618
rect 495234 640894 495854 665600
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 631820 495854 640338
rect 498954 644614 499574 665600
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 631820 499574 644058
rect 505794 651454 506414 665600
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 631820 506414 650898
rect 509514 655174 510134 665600
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 631820 510134 654618
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 631820 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 631820 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 631820 524414 632898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 631820 528134 636618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 478956 615454 479276 615486
rect 478956 615218 478998 615454
rect 479234 615218 479276 615454
rect 478956 615134 479276 615218
rect 478956 614898 478998 615134
rect 479234 614898 479276 615134
rect 478956 614866 479276 614898
rect 509676 615454 509996 615486
rect 509676 615218 509718 615454
rect 509954 615218 509996 615454
rect 509676 615134 509996 615218
rect 509676 614898 509718 615134
rect 509954 614898 509996 615134
rect 509676 614866 509996 614898
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 494316 597454 494636 597486
rect 494316 597218 494358 597454
rect 494594 597218 494636 597454
rect 494316 597134 494636 597218
rect 494316 596898 494358 597134
rect 494594 596898 494636 597134
rect 494316 596866 494636 596898
rect 525036 597454 525356 597486
rect 525036 597218 525078 597454
rect 525314 597218 525356 597454
rect 525036 597134 525356 597218
rect 525036 596898 525078 597134
rect 525314 596898 525356 597134
rect 525036 596866 525356 596898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 478956 579454 479276 579486
rect 478956 579218 478998 579454
rect 479234 579218 479276 579454
rect 478956 579134 479276 579218
rect 478956 578898 478998 579134
rect 479234 578898 479276 579134
rect 478956 578866 479276 578898
rect 509676 579454 509996 579486
rect 509676 579218 509718 579454
rect 509954 579218 509996 579454
rect 509676 579134 509996 579218
rect 509676 578898 509718 579134
rect 509954 578898 509996 579134
rect 509676 578866 509996 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 400000 470414 434898
rect 473514 547174 474134 573820
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 400000 474134 402618
rect 477234 550894 477854 573820
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 400000 477854 406338
rect 480954 554614 481574 573820
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 400000 481574 410058
rect 487794 561454 488414 573820
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 359568 381454 359888 381486
rect 359568 381218 359610 381454
rect 359846 381218 359888 381454
rect 359568 381134 359888 381218
rect 359568 380898 359610 381134
rect 359846 380898 359888 381134
rect 359568 380866 359888 380898
rect 390288 381454 390608 381486
rect 390288 381218 390330 381454
rect 390566 381218 390608 381454
rect 390288 381134 390608 381218
rect 390288 380898 390330 381134
rect 390566 380898 390608 381134
rect 390288 380866 390608 380898
rect 421008 381454 421328 381486
rect 421008 381218 421050 381454
rect 421286 381218 421328 381454
rect 421008 381134 421328 381218
rect 421008 380898 421050 381134
rect 421286 380898 421328 381134
rect 421008 380866 421328 380898
rect 451728 381454 452048 381486
rect 451728 381218 451770 381454
rect 452006 381218 452048 381454
rect 451728 381134 452048 381218
rect 451728 380898 451770 381134
rect 452006 380898 452048 381134
rect 451728 380866 452048 380898
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 344208 363454 344528 363486
rect 344208 363218 344250 363454
rect 344486 363218 344528 363454
rect 344208 363134 344528 363218
rect 344208 362898 344250 363134
rect 344486 362898 344528 363134
rect 344208 362866 344528 362898
rect 374928 363454 375248 363486
rect 374928 363218 374970 363454
rect 375206 363218 375248 363454
rect 374928 363134 375248 363218
rect 374928 362898 374970 363134
rect 375206 362898 375248 363134
rect 374928 362866 375248 362898
rect 405648 363454 405968 363486
rect 405648 363218 405690 363454
rect 405926 363218 405968 363454
rect 405648 363134 405968 363218
rect 405648 362898 405690 363134
rect 405926 362898 405968 363134
rect 405648 362866 405968 362898
rect 436368 363454 436688 363486
rect 436368 363218 436410 363454
rect 436646 363218 436688 363454
rect 436368 363134 436688 363218
rect 436368 362898 436410 363134
rect 436646 362898 436688 363134
rect 436368 362866 436688 362898
rect 467088 363454 467408 363486
rect 467088 363218 467130 363454
rect 467366 363218 467408 363454
rect 467088 363134 467408 363218
rect 467088 362898 467130 363134
rect 467366 362898 467408 363134
rect 467088 362866 467408 362898
rect 359568 345454 359888 345486
rect 359568 345218 359610 345454
rect 359846 345218 359888 345454
rect 359568 345134 359888 345218
rect 359568 344898 359610 345134
rect 359846 344898 359888 345134
rect 359568 344866 359888 344898
rect 390288 345454 390608 345486
rect 390288 345218 390330 345454
rect 390566 345218 390608 345454
rect 390288 345134 390608 345218
rect 390288 344898 390330 345134
rect 390566 344898 390608 345134
rect 390288 344866 390608 344898
rect 421008 345454 421328 345486
rect 421008 345218 421050 345454
rect 421286 345218 421328 345454
rect 421008 345134 421328 345218
rect 421008 344898 421050 345134
rect 421286 344898 421328 345134
rect 421008 344866 421328 344898
rect 451728 345454 452048 345486
rect 451728 345218 451770 345454
rect 452006 345218 452048 345454
rect 451728 345134 452048 345218
rect 451728 344898 451770 345134
rect 452006 344898 452048 345134
rect 451728 344866 452048 344898
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 344208 327454 344528 327486
rect 344208 327218 344250 327454
rect 344486 327218 344528 327454
rect 344208 327134 344528 327218
rect 344208 326898 344250 327134
rect 344486 326898 344528 327134
rect 344208 326866 344528 326898
rect 374928 327454 375248 327486
rect 374928 327218 374970 327454
rect 375206 327218 375248 327454
rect 374928 327134 375248 327218
rect 374928 326898 374970 327134
rect 375206 326898 375248 327134
rect 374928 326866 375248 326898
rect 405648 327454 405968 327486
rect 405648 327218 405690 327454
rect 405926 327218 405968 327454
rect 405648 327134 405968 327218
rect 405648 326898 405690 327134
rect 405926 326898 405968 327134
rect 405648 326866 405968 326898
rect 436368 327454 436688 327486
rect 436368 327218 436410 327454
rect 436646 327218 436688 327454
rect 436368 327134 436688 327218
rect 436368 326898 436410 327134
rect 436646 326898 436688 327134
rect 436368 326866 436688 326898
rect 467088 327454 467408 327486
rect 467088 327218 467130 327454
rect 467366 327218 467408 327454
rect 467088 327134 467408 327218
rect 467088 326898 467130 327134
rect 467366 326898 467408 327134
rect 467088 326866 467408 326898
rect 359568 309454 359888 309486
rect 359568 309218 359610 309454
rect 359846 309218 359888 309454
rect 359568 309134 359888 309218
rect 359568 308898 359610 309134
rect 359846 308898 359888 309134
rect 359568 308866 359888 308898
rect 390288 309454 390608 309486
rect 390288 309218 390330 309454
rect 390566 309218 390608 309454
rect 390288 309134 390608 309218
rect 390288 308898 390330 309134
rect 390566 308898 390608 309134
rect 390288 308866 390608 308898
rect 421008 309454 421328 309486
rect 421008 309218 421050 309454
rect 421286 309218 421328 309454
rect 421008 309134 421328 309218
rect 421008 308898 421050 309134
rect 421286 308898 421328 309134
rect 421008 308866 421328 308898
rect 451728 309454 452048 309486
rect 451728 309218 451770 309454
rect 452006 309218 452048 309454
rect 451728 309134 452048 309218
rect 451728 308898 451770 309134
rect 452006 308898 452048 309134
rect 451728 308866 452048 308898
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 344208 291454 344528 291486
rect 344208 291218 344250 291454
rect 344486 291218 344528 291454
rect 344208 291134 344528 291218
rect 344208 290898 344250 291134
rect 344486 290898 344528 291134
rect 344208 290866 344528 290898
rect 374928 291454 375248 291486
rect 374928 291218 374970 291454
rect 375206 291218 375248 291454
rect 374928 291134 375248 291218
rect 374928 290898 374970 291134
rect 375206 290898 375248 291134
rect 374928 290866 375248 290898
rect 405648 291454 405968 291486
rect 405648 291218 405690 291454
rect 405926 291218 405968 291454
rect 405648 291134 405968 291218
rect 405648 290898 405690 291134
rect 405926 290898 405968 291134
rect 405648 290866 405968 290898
rect 436368 291454 436688 291486
rect 436368 291218 436410 291454
rect 436646 291218 436688 291454
rect 436368 291134 436688 291218
rect 436368 290898 436410 291134
rect 436646 290898 436688 291134
rect 436368 290866 436688 290898
rect 467088 291454 467408 291486
rect 467088 291218 467130 291454
rect 467366 291218 467408 291454
rect 467088 291134 467408 291218
rect 467088 290898 467130 291134
rect 467366 290898 467408 291134
rect 467088 290866 467408 290898
rect 359568 273454 359888 273486
rect 359568 273218 359610 273454
rect 359846 273218 359888 273454
rect 359568 273134 359888 273218
rect 359568 272898 359610 273134
rect 359846 272898 359888 273134
rect 359568 272866 359888 272898
rect 390288 273454 390608 273486
rect 390288 273218 390330 273454
rect 390566 273218 390608 273454
rect 390288 273134 390608 273218
rect 390288 272898 390330 273134
rect 390566 272898 390608 273134
rect 390288 272866 390608 272898
rect 421008 273454 421328 273486
rect 421008 273218 421050 273454
rect 421286 273218 421328 273454
rect 421008 273134 421328 273218
rect 421008 272898 421050 273134
rect 421286 272898 421328 273134
rect 421008 272866 421328 272898
rect 451728 273454 452048 273486
rect 451728 273218 451770 273454
rect 452006 273218 452048 273454
rect 451728 273134 452048 273218
rect 451728 272898 451770 273134
rect 452006 272898 452048 273134
rect 451728 272866 452048 272898
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 237454 344414 256000
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 241174 348134 256000
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 244894 351854 256000
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 248614 355574 256000
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 255454 362414 256000
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 223174 366134 256000
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 226894 369854 256000
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 230614 373574 256000
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 237454 380414 256000
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 241174 384134 256000
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 244894 387854 256000
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 248614 391574 256000
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 255454 398414 256000
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 223174 402134 256000
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 226894 405854 256000
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 230614 409574 256000
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 237454 416414 256000
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 241174 420134 256000
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 244894 423854 256000
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 248614 427574 256000
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 255454 434414 256000
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 223174 438134 256000
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 226894 441854 256000
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 230614 445574 256000
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 237454 452414 256000
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 241174 456134 256000
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 244894 459854 256000
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 248614 463574 256000
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 255454 470414 256000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 461648 223174 461968 223206
rect 461648 222938 461690 223174
rect 461926 222938 461968 223174
rect 461648 222854 461968 222938
rect 461648 222618 461690 222854
rect 461926 222618 461968 222854
rect 461648 222586 461968 222618
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 461648 187174 461968 187206
rect 461648 186938 461690 187174
rect 461926 186938 461968 187174
rect 461648 186854 461968 186938
rect 461648 186618 461690 186854
rect 461926 186618 461968 186854
rect 461648 186586 461968 186618
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 461648 151174 461968 151206
rect 461648 150938 461690 151174
rect 461926 150938 461968 151174
rect 461648 150854 461968 150938
rect 461648 150618 461690 150854
rect 461926 150618 461968 150854
rect 461648 150586 461968 150618
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 461648 115174 461968 115206
rect 461648 114938 461690 115174
rect 461926 114938 461968 115174
rect 461648 114854 461968 114938
rect 461648 114618 461690 114854
rect 461926 114618 461968 114854
rect 461648 114586 461968 114618
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 461648 79174 461968 79206
rect 461648 78938 461690 79174
rect 461926 78938 461968 79174
rect 461648 78854 461968 78938
rect 461648 78618 461690 78854
rect 461926 78618 461968 78854
rect 461648 78586 461968 78618
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 461648 43174 461968 43206
rect 461648 42938 461690 43174
rect 461926 42938 461968 43174
rect 461648 42854 461968 42938
rect 461648 42618 461690 42854
rect 461926 42618 461968 42854
rect 461648 42586 461968 42618
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 458403 3364 458469 3365
rect 458403 3300 458404 3364
rect 458468 3300 458469 3364
rect 458403 3299 458469 3300
rect 458406 2957 458466 3299
rect 458403 2956 458469 2957
rect 458403 2892 458404 2956
rect 458468 2892 458469 2956
rect 458403 2891 458469 2892
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 -7066 460454 28938
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 461648 7174 461968 7206
rect 461648 6938 461690 7174
rect 461926 6938 461968 7174
rect 461648 6854 461968 6938
rect 461648 6618 461690 6854
rect 461926 6618 461968 6854
rect 461648 6586 461968 6618
rect 462635 3636 462701 3637
rect 462635 3572 462636 3636
rect 462700 3572 462701 3636
rect 462635 3571 462701 3572
rect 462638 2685 462698 3571
rect 463739 3500 463805 3501
rect 463739 3436 463740 3500
rect 463804 3436 463805 3500
rect 463739 3435 463805 3436
rect 469794 3454 470414 38898
rect 463742 2821 463802 3435
rect 467235 3364 467301 3365
rect 467235 3300 467236 3364
rect 467300 3300 467301 3364
rect 467235 3299 467301 3300
rect 466315 3228 466381 3229
rect 466315 3164 466316 3228
rect 466380 3164 466381 3228
rect 466315 3163 466381 3164
rect 463739 2820 463805 2821
rect 463739 2756 463740 2820
rect 463804 2756 463805 2820
rect 463739 2755 463805 2756
rect 462635 2684 462701 2685
rect 462635 2620 462636 2684
rect 462700 2620 462701 2684
rect 462635 2619 462701 2620
rect 466318 2549 466378 3163
rect 467238 2549 467298 3299
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 466315 2548 466381 2549
rect 466315 2484 466316 2548
rect 466380 2484 466381 2548
rect 466315 2483 466381 2484
rect 467235 2548 467301 2549
rect 467235 2484 467236 2548
rect 467300 2484 467301 2548
rect 467235 2483 467301 2484
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 223174 474134 256000
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 226894 477854 256000
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 230614 481574 256000
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 565174 492134 573820
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 568894 495854 573820
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 572614 499574 573820
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 543454 506414 573820
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 547174 510134 573820
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 498147 3092 498213 3093
rect 498147 3028 498148 3092
rect 498212 3028 498213 3092
rect 498147 3027 498213 3028
rect 498150 2549 498210 3027
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 498147 2548 498213 2549
rect 498147 2484 498148 2548
rect 498212 2484 498213 2548
rect 498147 2483 498213 2484
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 550894 513854 573820
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 554614 517574 573820
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 561454 524414 573820
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 565174 528134 573820
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 538448 327454 538768 327486
rect 538448 327218 538490 327454
rect 538726 327218 538768 327454
rect 538448 327134 538768 327218
rect 538448 326898 538490 327134
rect 538726 326898 538768 327134
rect 538448 326866 538768 326898
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 538448 291454 538768 291486
rect 538448 291218 538490 291454
rect 538726 291218 538768 291454
rect 538448 291134 538768 291218
rect 538448 290898 538490 291134
rect 538726 290898 538768 291134
rect 538448 290866 538768 290898
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 538448 255454 538768 255486
rect 538448 255218 538490 255454
rect 538726 255218 538768 255454
rect 538448 255134 538768 255218
rect 538448 254898 538490 255134
rect 538726 254898 538768 255134
rect 538448 254866 538768 254898
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 538448 219454 538768 219486
rect 538448 219218 538490 219454
rect 538726 219218 538768 219454
rect 538448 219134 538768 219218
rect 538448 218898 538490 219134
rect 538726 218898 538768 219134
rect 538448 218866 538768 218898
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 538448 183454 538768 183486
rect 538448 183218 538490 183454
rect 538726 183218 538768 183454
rect 538448 183134 538768 183218
rect 538448 182898 538490 183134
rect 538726 182898 538768 183134
rect 538448 182866 538768 182898
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 538448 147454 538768 147486
rect 538448 147218 538490 147454
rect 538726 147218 538768 147454
rect 538448 147134 538768 147218
rect 538448 146898 538490 147134
rect 538726 146898 538768 147134
rect 538448 146866 538768 146898
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 538448 111454 538768 111486
rect 538448 111218 538490 111454
rect 538726 111218 538768 111454
rect 538448 111134 538768 111218
rect 538448 110898 538490 111134
rect 538726 110898 538768 111134
rect 538448 110866 538768 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 538448 75454 538768 75486
rect 538448 75218 538490 75454
rect 538726 75218 538768 75454
rect 538448 75134 538768 75218
rect 538448 74898 538490 75134
rect 538726 74898 538768 75134
rect 538448 74866 538768 74898
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 538448 39454 538768 39486
rect 538448 39218 538490 39454
rect 538726 39218 538768 39454
rect 538448 39134 538768 39218
rect 538448 38898 538490 39134
rect 538726 38898 538768 39134
rect 538448 38866 538768 38898
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 529979 3228 530045 3229
rect 529979 3164 529980 3228
rect 530044 3164 530045 3228
rect 529979 3163 530045 3164
rect 529982 2685 530042 3163
rect 529979 2684 530045 2685
rect 529979 2620 529980 2684
rect 530044 2620 530045 2684
rect 529979 2619 530045 2620
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 -7066 532454 28938
rect 533475 3772 533541 3773
rect 533475 3708 533476 3772
rect 533540 3708 533541 3772
rect 533475 3707 533541 3708
rect 533478 2957 533538 3707
rect 541794 3454 542414 38898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545251 3636 545317 3637
rect 545251 3572 545252 3636
rect 545316 3572 545317 3636
rect 545251 3571 545317 3572
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 533475 2956 533541 2957
rect 533475 2892 533476 2956
rect 533540 2892 533541 2956
rect 533475 2891 533541 2892
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 533291 2820 533357 2821
rect 533291 2756 533292 2820
rect 533356 2756 533357 2820
rect 533291 2755 533357 2756
rect 533294 2685 533354 2755
rect 533291 2684 533357 2685
rect 533291 2620 533292 2684
rect 533356 2620 533357 2684
rect 533291 2619 533357 2620
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 -346 542414 2898
rect 545254 2549 545314 3571
rect 545251 2548 545317 2549
rect 545251 2484 545252 2548
rect 545316 2484 545317 2548
rect 545251 2483 545317 2484
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 -1306 546134 6618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 547643 3500 547709 3501
rect 547643 3436 547644 3500
rect 547708 3436 547709 3500
rect 547643 3435 547709 3436
rect 547646 2549 547706 3435
rect 547643 2548 547709 2549
rect 547643 2484 547644 2548
rect 547708 2484 547709 2548
rect 547643 2483 547709 2484
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 -2266 549854 10338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 553808 331174 554128 331206
rect 553808 330938 553850 331174
rect 554086 330938 554128 331174
rect 553808 330854 554128 330938
rect 553808 330618 553850 330854
rect 554086 330618 554128 330854
rect 553808 330586 554128 330618
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 553808 295174 554128 295206
rect 553808 294938 553850 295174
rect 554086 294938 554128 295174
rect 553808 294854 554128 294938
rect 553808 294618 553850 294854
rect 554086 294618 554128 294854
rect 553808 294586 554128 294618
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 553808 259174 554128 259206
rect 553808 258938 553850 259174
rect 554086 258938 554128 259174
rect 553808 258854 554128 258938
rect 553808 258618 553850 258854
rect 554086 258618 554128 258854
rect 553808 258586 554128 258618
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 553808 223174 554128 223206
rect 553808 222938 553850 223174
rect 554086 222938 554128 223174
rect 553808 222854 554128 222938
rect 553808 222618 553850 222854
rect 554086 222618 554128 222854
rect 553808 222586 554128 222618
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 553808 187174 554128 187206
rect 553808 186938 553850 187174
rect 554086 186938 554128 187174
rect 553808 186854 554128 186938
rect 553808 186618 553850 186854
rect 554086 186618 554128 186854
rect 553808 186586 554128 186618
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 553808 151174 554128 151206
rect 553808 150938 553850 151174
rect 554086 150938 554128 151174
rect 553808 150854 554128 150938
rect 553808 150618 553850 150854
rect 554086 150618 554128 150854
rect 553808 150586 554128 150618
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 553808 115174 554128 115206
rect 553808 114938 553850 115174
rect 554086 114938 554128 115174
rect 553808 114854 554128 114938
rect 553808 114618 553850 114854
rect 554086 114618 554128 114854
rect 553808 114586 554128 114618
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 553808 79174 554128 79206
rect 553808 78938 553850 79174
rect 554086 78938 554128 79174
rect 553808 78854 554128 78938
rect 553808 78618 553850 78854
rect 554086 78618 554128 78854
rect 553808 78586 554128 78618
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 553808 43174 554128 43206
rect 553808 42938 553850 43174
rect 554086 42938 554128 43174
rect 553808 42854 554128 42938
rect 553808 42618 553850 42854
rect 554086 42618 554128 42854
rect 553808 42586 554128 42618
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552427 3364 552493 3365
rect 552427 3300 552428 3364
rect 552492 3300 552493 3364
rect 552427 3299 552493 3300
rect 552430 2685 552490 3299
rect 552427 2684 552493 2685
rect 552427 2620 552428 2684
rect 552492 2620 552493 2684
rect 552427 2619 552493 2620
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 -3226 553574 14058
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 553808 7174 554128 7206
rect 553808 6938 553850 7174
rect 554086 6938 554128 7174
rect 553808 6854 554128 6938
rect 553808 6618 553850 6854
rect 554086 6618 554128 6854
rect 553808 6586 554128 6618
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 -4186 557294 17778
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 558499 3908 558565 3909
rect 558499 3844 558500 3908
rect 558564 3844 558565 3908
rect 558499 3843 558565 3844
rect 558502 2821 558562 3843
rect 558499 2820 558565 2821
rect 558499 2756 558500 2820
rect 558564 2756 558565 2820
rect 558499 2755 558565 2756
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 574691 344724 574757 344725
rect 574691 344660 574692 344724
rect 574756 344660 574757 344724
rect 574691 344659 574757 344660
rect 569168 327454 569488 327486
rect 569168 327218 569210 327454
rect 569446 327218 569488 327454
rect 569168 327134 569488 327218
rect 569168 326898 569210 327134
rect 569446 326898 569488 327134
rect 569168 326866 569488 326898
rect 574694 325277 574754 344659
rect 574875 330308 574941 330309
rect 574875 330244 574876 330308
rect 574940 330244 574941 330308
rect 574875 330243 574941 330244
rect 574691 325276 574757 325277
rect 574691 325212 574692 325276
rect 574756 325212 574757 325276
rect 574691 325211 574757 325212
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 574878 312085 574938 330243
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 575059 315892 575125 315893
rect 575059 315828 575060 315892
rect 575124 315828 575125 315892
rect 575059 315827 575125 315828
rect 574875 312084 574941 312085
rect 574875 312020 574876 312084
rect 574940 312020 574941 312084
rect 574875 312019 574941 312020
rect 574691 301476 574757 301477
rect 574691 301412 574692 301476
rect 574756 301412 574757 301476
rect 574691 301411 574757 301412
rect 569168 291454 569488 291486
rect 569168 291218 569210 291454
rect 569446 291218 569488 291454
rect 569168 291134 569488 291218
rect 569168 290898 569210 291134
rect 569446 290898 569488 291134
rect 569168 290866 569488 290898
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 574694 272237 574754 301411
rect 575062 298757 575122 315827
rect 575059 298756 575125 298757
rect 575059 298692 575060 298756
rect 575124 298692 575125 298756
rect 575059 298691 575125 298692
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 575059 287060 575125 287061
rect 575059 286996 575060 287060
rect 575124 286996 575125 287060
rect 575059 286995 575125 286996
rect 574875 272644 574941 272645
rect 574875 272580 574876 272644
rect 574940 272580 574941 272644
rect 574875 272579 574941 272580
rect 574691 272236 574757 272237
rect 574691 272172 574692 272236
rect 574756 272172 574757 272236
rect 574691 272171 574757 272172
rect 574691 258228 574757 258229
rect 574691 258164 574692 258228
rect 574756 258164 574757 258228
rect 574691 258163 574757 258164
rect 569168 255454 569488 255486
rect 569168 255218 569210 255454
rect 569446 255218 569488 255454
rect 569168 255134 569488 255218
rect 569168 254898 569210 255134
rect 569446 254898 569488 255134
rect 569168 254866 569488 254898
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 574694 232389 574754 258163
rect 574878 245581 574938 272579
rect 575062 258909 575122 286995
rect 575059 258908 575125 258909
rect 575059 258844 575060 258908
rect 575124 258844 575125 258908
rect 575059 258843 575125 258844
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 574875 245580 574941 245581
rect 574875 245516 574876 245580
rect 574940 245516 574941 245580
rect 574875 245515 574941 245516
rect 574875 243812 574941 243813
rect 574875 243748 574876 243812
rect 574940 243748 574941 243812
rect 574875 243747 574941 243748
rect 574691 232388 574757 232389
rect 574691 232324 574692 232388
rect 574756 232324 574757 232388
rect 574691 232323 574757 232324
rect 574691 229396 574757 229397
rect 574691 229332 574692 229396
rect 574756 229332 574757 229396
rect 574691 229331 574757 229332
rect 569168 219454 569488 219486
rect 569168 219218 569210 219454
rect 569446 219218 569488 219454
rect 569168 219134 569488 219218
rect 569168 218898 569210 219134
rect 569446 218898 569488 219134
rect 569168 218866 569488 218898
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 574694 205733 574754 229331
rect 574878 219061 574938 243747
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 574875 219060 574941 219061
rect 574875 218996 574876 219060
rect 574940 218996 574941 219060
rect 574875 218995 574941 218996
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 574875 214980 574941 214981
rect 574875 214916 574876 214980
rect 574940 214916 574941 214980
rect 574875 214915 574941 214916
rect 574691 205732 574757 205733
rect 574691 205668 574692 205732
rect 574756 205668 574757 205732
rect 574691 205667 574757 205668
rect 574691 200564 574757 200565
rect 574691 200500 574692 200564
rect 574756 200500 574757 200564
rect 574691 200499 574757 200500
rect 569168 183454 569488 183486
rect 569168 183218 569210 183454
rect 569446 183218 569488 183454
rect 569168 183134 569488 183218
rect 569168 182898 569210 183134
rect 569446 182898 569488 183134
rect 569168 182866 569488 182898
rect 574694 179213 574754 200499
rect 574878 192541 574938 214915
rect 574875 192540 574941 192541
rect 574875 192476 574876 192540
rect 574940 192476 574941 192540
rect 574875 192475 574941 192476
rect 574875 186148 574941 186149
rect 574875 186084 574876 186148
rect 574940 186084 574941 186148
rect 574875 186083 574941 186084
rect 574691 179212 574757 179213
rect 574691 179148 574692 179212
rect 574756 179148 574757 179212
rect 574691 179147 574757 179148
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 574691 171732 574757 171733
rect 574691 171668 574692 171732
rect 574756 171668 574757 171732
rect 574691 171667 574757 171668
rect 574694 152693 574754 171667
rect 574878 165885 574938 186083
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 574875 165884 574941 165885
rect 574875 165820 574876 165884
rect 574940 165820 574941 165884
rect 574875 165819 574941 165820
rect 574875 157316 574941 157317
rect 574875 157252 574876 157316
rect 574940 157252 574941 157316
rect 574875 157251 574941 157252
rect 574691 152692 574757 152693
rect 574691 152628 574692 152692
rect 574756 152628 574757 152692
rect 574691 152627 574757 152628
rect 569168 147454 569488 147486
rect 569168 147218 569210 147454
rect 569446 147218 569488 147454
rect 569168 147134 569488 147218
rect 569168 146898 569210 147134
rect 569446 146898 569488 147134
rect 569168 146866 569488 146898
rect 574691 142900 574757 142901
rect 574691 142836 574692 142900
rect 574756 142836 574757 142900
rect 574691 142835 574757 142836
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 574694 126037 574754 142835
rect 574878 139365 574938 157251
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 574875 139364 574941 139365
rect 574875 139300 574876 139364
rect 574940 139300 574941 139364
rect 574875 139299 574941 139300
rect 574875 128484 574941 128485
rect 574875 128420 574876 128484
rect 574940 128420 574941 128484
rect 574875 128419 574941 128420
rect 574691 126036 574757 126037
rect 574691 125972 574692 126036
rect 574756 125972 574757 126036
rect 574691 125971 574757 125972
rect 574691 114068 574757 114069
rect 574691 114004 574692 114068
rect 574756 114004 574757 114068
rect 574691 114003 574757 114004
rect 569168 111454 569488 111486
rect 569168 111218 569210 111454
rect 569446 111218 569488 111454
rect 569168 111134 569488 111218
rect 569168 110898 569210 111134
rect 569446 110898 569488 111134
rect 569168 110866 569488 110898
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 574694 99517 574754 114003
rect 574878 112845 574938 128419
rect 574875 112844 574941 112845
rect 574875 112780 574876 112844
rect 574940 112780 574941 112844
rect 574875 112779 574941 112780
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 574875 99652 574941 99653
rect 574875 99588 574876 99652
rect 574940 99588 574941 99652
rect 574875 99587 574941 99588
rect 574691 99516 574757 99517
rect 574691 99452 574692 99516
rect 574756 99452 574757 99516
rect 574691 99451 574757 99452
rect 574878 86189 574938 99587
rect 574875 86188 574941 86189
rect 574875 86124 574876 86188
rect 574940 86124 574941 86188
rect 574875 86123 574941 86124
rect 574691 85236 574757 85237
rect 574691 85172 574692 85236
rect 574756 85172 574757 85236
rect 574691 85171 574757 85172
rect 569168 75454 569488 75486
rect 569168 75218 569210 75454
rect 569446 75218 569488 75454
rect 569168 75134 569488 75218
rect 569168 74898 569210 75134
rect 569446 74898 569488 75134
rect 569168 74866 569488 74898
rect 574694 72997 574754 85171
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 574691 72996 574757 72997
rect 574691 72932 574692 72996
rect 574756 72932 574757 72996
rect 574691 72931 574757 72932
rect 574691 70820 574757 70821
rect 574691 70756 574692 70820
rect 574756 70756 574757 70820
rect 574691 70755 574757 70756
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 574694 59669 574754 70755
rect 574691 59668 574757 59669
rect 574691 59604 574692 59668
rect 574756 59604 574757 59668
rect 574691 59603 574757 59604
rect 574691 56404 574757 56405
rect 574691 56340 574692 56404
rect 574756 56340 574757 56404
rect 574691 56339 574757 56340
rect 574694 46341 574754 56339
rect 574691 46340 574757 46341
rect 574691 46276 574692 46340
rect 574756 46276 574757 46340
rect 574691 46275 574757 46276
rect 574691 41988 574757 41989
rect 574691 41924 574692 41988
rect 574756 41924 574757 41988
rect 574691 41923 574757 41924
rect 569168 39454 569488 39486
rect 569168 39218 569210 39454
rect 569446 39218 569488 39454
rect 569168 39134 569488 39218
rect 569168 38898 569210 39134
rect 569446 38898 569488 39134
rect 569168 38866 569488 38898
rect 574694 33149 574754 41923
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 574691 33148 574757 33149
rect 574691 33084 574692 33148
rect 574756 33084 574757 33148
rect 574691 33083 574757 33084
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 575427 27572 575493 27573
rect 575427 27508 575428 27572
rect 575492 27508 575493 27572
rect 575427 27507 575493 27508
rect 575430 19821 575490 27507
rect 575427 19820 575493 19821
rect 575427 19756 575428 19820
rect 575492 19756 575493 19820
rect 575427 19755 575493 19756
rect 574691 13156 574757 13157
rect 574691 13092 574692 13156
rect 574756 13092 574757 13156
rect 574691 13091 574757 13092
rect 574694 6629 574754 13091
rect 574691 6628 574757 6629
rect 574691 6564 574692 6628
rect 574756 6564 574757 6628
rect 574691 6563 574757 6564
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 85922 687218 86158 687454
rect 85922 686898 86158 687134
rect 88522 687218 88758 687454
rect 88522 686898 88758 687134
rect 95722 687218 95958 687454
rect 95722 686898 95958 687134
rect 102922 687218 103158 687454
rect 102922 686898 103158 687134
rect 110122 687218 110358 687454
rect 110122 686898 110358 687134
rect 117322 687218 117558 687454
rect 117322 686898 117558 687134
rect 119922 687218 120158 687454
rect 119922 686898 120158 687134
rect 84922 669218 85158 669454
rect 84922 668898 85158 669134
rect 92122 669218 92358 669454
rect 92122 668898 92358 669134
rect 99322 669218 99558 669454
rect 99322 668898 99558 669134
rect 106522 669218 106758 669454
rect 106522 668898 106758 669134
rect 113722 669218 113958 669454
rect 113722 668898 113958 669134
rect 120922 669218 121158 669454
rect 120922 668898 121158 669134
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 79542 615218 79778 615454
rect 79542 614898 79778 615134
rect 110262 615218 110498 615454
rect 110262 614898 110498 615134
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 94902 597218 95138 597454
rect 94902 596898 95138 597134
rect 125622 597218 125858 597454
rect 125622 596898 125858 597134
rect 79542 579218 79778 579454
rect 79542 578898 79778 579134
rect 110262 579218 110498 579454
rect 110262 578898 110498 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 21008 399218 21244 399454
rect 21008 398898 21244 399134
rect 155376 399218 155612 399454
rect 155376 398898 155612 399134
rect 20328 381218 20564 381454
rect 20328 380898 20564 381134
rect 156056 381218 156292 381454
rect 156056 380898 156292 381134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 21008 363218 21244 363454
rect 21008 362898 21244 363134
rect 155376 363218 155612 363454
rect 155376 362898 155612 363134
rect 20328 345218 20564 345454
rect 20328 344898 20564 345134
rect 156056 345218 156292 345454
rect 156056 344898 156292 345134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 21008 327218 21244 327454
rect 21008 326898 21244 327134
rect 155376 327218 155612 327454
rect 155376 326898 155612 327134
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 30986 301438 31222 301674
rect 31306 301438 31542 301674
rect 30986 301118 31222 301354
rect 31306 301118 31542 301354
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 301438 67222 301674
rect 67306 301438 67542 301674
rect 66986 301118 67222 301354
rect 67306 301118 67542 301354
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 301438 103222 301674
rect 103306 301438 103542 301674
rect 102986 301118 103222 301354
rect 103306 301118 103542 301354
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 138986 301438 139222 301674
rect 139306 301438 139542 301674
rect 138986 301118 139222 301354
rect 139306 301118 139542 301354
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 20328 273218 20564 273454
rect 20328 272898 20564 273134
rect 156056 273218 156292 273454
rect 156056 272898 156292 273134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 21008 255218 21244 255454
rect 21008 254898 21244 255134
rect 155376 255218 155612 255454
rect 155376 254898 155612 255134
rect 20328 237218 20564 237454
rect 20328 236898 20564 237134
rect 156056 237218 156292 237454
rect 156056 236898 156292 237134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 21008 219218 21244 219454
rect 21008 218898 21244 219134
rect 155376 219218 155612 219454
rect 155376 218898 155612 219134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 241162 687218 241398 687454
rect 241162 686898 241398 687134
rect 243762 687218 243998 687454
rect 243762 686898 243998 687134
rect 250962 687218 251198 687454
rect 250962 686898 251198 687134
rect 258162 687218 258398 687454
rect 258162 686898 258398 687134
rect 265362 687218 265598 687454
rect 265362 686898 265598 687134
rect 272562 687218 272798 687454
rect 272562 686898 272798 687134
rect 275162 687218 275398 687454
rect 275162 686898 275398 687134
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 240162 669218 240398 669454
rect 240162 668898 240398 669134
rect 247362 669218 247598 669454
rect 247362 668898 247598 669134
rect 254562 669218 254798 669454
rect 254562 668898 254798 669134
rect 261762 669218 261998 669454
rect 261762 668898 261998 669134
rect 268962 669218 269198 669454
rect 268962 668898 269198 669134
rect 276162 669218 276398 669454
rect 276162 668898 276398 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 239450 615218 239686 615454
rect 239450 614898 239686 615134
rect 270170 615218 270406 615454
rect 270170 614898 270406 615134
rect 254810 597218 255046 597454
rect 254810 596898 255046 597134
rect 285530 597218 285766 597454
rect 285530 596898 285766 597134
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 239450 579218 239686 579454
rect 239450 578898 239686 579134
rect 270170 579218 270406 579454
rect 270170 578898 270406 579134
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 181008 399218 181244 399454
rect 181008 398898 181244 399134
rect 315376 399218 315612 399454
rect 315376 398898 315612 399134
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 180328 381218 180564 381454
rect 180328 380898 180564 381134
rect 316056 381218 316292 381454
rect 316056 380898 316292 381134
rect 181008 363218 181244 363454
rect 181008 362898 181244 363134
rect 315376 363218 315612 363454
rect 315376 362898 315612 363134
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 180328 345218 180564 345454
rect 180328 344898 180564 345134
rect 316056 345218 316292 345454
rect 316056 344898 316292 345134
rect 181008 327218 181244 327454
rect 181008 326898 181244 327134
rect 315376 327218 315612 327454
rect 315376 326898 315612 327134
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 301438 175222 301674
rect 175306 301438 175542 301674
rect 174986 301118 175222 301354
rect 175306 301118 175542 301354
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 301438 211222 301674
rect 211306 301438 211542 301674
rect 210986 301118 211222 301354
rect 211306 301118 211542 301354
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 301438 247222 301674
rect 247306 301438 247542 301674
rect 246986 301118 247222 301354
rect 247306 301118 247542 301354
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 282986 301438 283222 301674
rect 283306 301438 283542 301674
rect 282986 301118 283222 301354
rect 283306 301118 283542 301354
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 180328 273218 180564 273454
rect 180328 272898 180564 273134
rect 316056 273218 316292 273454
rect 316056 272898 316292 273134
rect 181008 255218 181244 255454
rect 181008 254898 181244 255134
rect 315376 255218 315612 255454
rect 315376 254898 315612 255134
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 180328 237218 180564 237454
rect 180328 236898 180564 237134
rect 316056 237218 316292 237454
rect 316056 236898 316292 237134
rect 181008 219218 181244 219454
rect 181008 218898 181244 219134
rect 315376 219218 315612 219454
rect 315376 218898 315612 219134
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 486322 687218 486558 687454
rect 486322 686898 486558 687134
rect 489922 687218 490158 687454
rect 489922 686898 490158 687134
rect 495522 687218 495758 687454
rect 495522 686898 495758 687134
rect 501122 687218 501358 687454
rect 501122 686898 501358 687134
rect 506722 687218 506958 687454
rect 506722 686898 506958 687134
rect 510322 687218 510558 687454
rect 510322 686898 510558 687134
rect 487122 669218 487358 669454
rect 487122 668898 487358 669134
rect 492722 669218 492958 669454
rect 492722 668898 492958 669134
rect 498322 669218 498558 669454
rect 498322 668898 498558 669134
rect 503922 669218 504158 669454
rect 503922 668898 504158 669134
rect 509522 669218 509758 669454
rect 509522 668898 509758 669134
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 478998 615218 479234 615454
rect 478998 614898 479234 615134
rect 509718 615218 509954 615454
rect 509718 614898 509954 615134
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 494358 597218 494594 597454
rect 494358 596898 494594 597134
rect 525078 597218 525314 597454
rect 525078 596898 525314 597134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 478998 579218 479234 579454
rect 478998 578898 479234 579134
rect 509718 579218 509954 579454
rect 509718 578898 509954 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 359610 381218 359846 381454
rect 359610 380898 359846 381134
rect 390330 381218 390566 381454
rect 390330 380898 390566 381134
rect 421050 381218 421286 381454
rect 421050 380898 421286 381134
rect 451770 381218 452006 381454
rect 451770 380898 452006 381134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 344250 363218 344486 363454
rect 344250 362898 344486 363134
rect 374970 363218 375206 363454
rect 374970 362898 375206 363134
rect 405690 363218 405926 363454
rect 405690 362898 405926 363134
rect 436410 363218 436646 363454
rect 436410 362898 436646 363134
rect 467130 363218 467366 363454
rect 467130 362898 467366 363134
rect 359610 345218 359846 345454
rect 359610 344898 359846 345134
rect 390330 345218 390566 345454
rect 390330 344898 390566 345134
rect 421050 345218 421286 345454
rect 421050 344898 421286 345134
rect 451770 345218 452006 345454
rect 451770 344898 452006 345134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 344250 327218 344486 327454
rect 344250 326898 344486 327134
rect 374970 327218 375206 327454
rect 374970 326898 375206 327134
rect 405690 327218 405926 327454
rect 405690 326898 405926 327134
rect 436410 327218 436646 327454
rect 436410 326898 436646 327134
rect 467130 327218 467366 327454
rect 467130 326898 467366 327134
rect 359610 309218 359846 309454
rect 359610 308898 359846 309134
rect 390330 309218 390566 309454
rect 390330 308898 390566 309134
rect 421050 309218 421286 309454
rect 421050 308898 421286 309134
rect 451770 309218 452006 309454
rect 451770 308898 452006 309134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 344250 291218 344486 291454
rect 344250 290898 344486 291134
rect 374970 291218 375206 291454
rect 374970 290898 375206 291134
rect 405690 291218 405926 291454
rect 405690 290898 405926 291134
rect 436410 291218 436646 291454
rect 436410 290898 436646 291134
rect 467130 291218 467366 291454
rect 467130 290898 467366 291134
rect 359610 273218 359846 273454
rect 359610 272898 359846 273134
rect 390330 273218 390566 273454
rect 390330 272898 390566 273134
rect 421050 273218 421286 273454
rect 421050 272898 421286 273134
rect 451770 273218 452006 273454
rect 451770 272898 452006 273134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 461690 222938 461926 223174
rect 461690 222618 461926 222854
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 461690 186938 461926 187174
rect 461690 186618 461926 186854
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 461690 150938 461926 151174
rect 461690 150618 461926 150854
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 461690 114938 461926 115174
rect 461690 114618 461926 114854
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 461690 78938 461926 79174
rect 461690 78618 461926 78854
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 461690 42938 461926 43174
rect 461690 42618 461926 42854
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 461690 6938 461926 7174
rect 461690 6618 461926 6854
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 538490 327218 538726 327454
rect 538490 326898 538726 327134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 538490 291218 538726 291454
rect 538490 290898 538726 291134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 538490 255218 538726 255454
rect 538490 254898 538726 255134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 538490 219218 538726 219454
rect 538490 218898 538726 219134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 538490 183218 538726 183454
rect 538490 182898 538726 183134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 538490 147218 538726 147454
rect 538490 146898 538726 147134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 538490 111218 538726 111454
rect 538490 110898 538726 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 538490 75218 538726 75454
rect 538490 74898 538726 75134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 538490 39218 538726 39454
rect 538490 38898 538726 39134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 553850 330938 554086 331174
rect 553850 330618 554086 330854
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 553850 294938 554086 295174
rect 553850 294618 554086 294854
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 553850 258938 554086 259174
rect 553850 258618 554086 258854
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 553850 222938 554086 223174
rect 553850 222618 554086 222854
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 553850 186938 554086 187174
rect 553850 186618 554086 186854
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 553850 150938 554086 151174
rect 553850 150618 554086 150854
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 553850 114938 554086 115174
rect 553850 114618 554086 114854
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 553850 78938 554086 79174
rect 553850 78618 554086 78854
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 553850 42938 554086 43174
rect 553850 42618 554086 42854
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 553850 6938 554086 7174
rect 553850 6618 554086 6854
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 569210 327218 569446 327454
rect 569210 326898 569446 327134
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 569210 291218 569446 291454
rect 569210 290898 569446 291134
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 569210 255218 569446 255454
rect 569210 254898 569446 255134
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 569210 219218 569446 219454
rect 569210 218898 569446 219134
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 569210 183218 569446 183454
rect 569210 182898 569446 183134
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 569210 147218 569446 147454
rect 569210 146898 569446 147134
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 569210 111218 569446 111454
rect 569210 110898 569446 111134
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 569210 75218 569446 75454
rect 569210 74898 569446 75134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 569210 39218 569446 39454
rect 569210 38898 569446 39134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 85922 687454
rect 86158 687218 88522 687454
rect 88758 687218 95722 687454
rect 95958 687218 102922 687454
rect 103158 687218 110122 687454
rect 110358 687218 117322 687454
rect 117558 687218 119922 687454
rect 120158 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 241162 687454
rect 241398 687218 243762 687454
rect 243998 687218 250962 687454
rect 251198 687218 258162 687454
rect 258398 687218 265362 687454
rect 265598 687218 272562 687454
rect 272798 687218 275162 687454
rect 275398 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 486322 687454
rect 486558 687218 489922 687454
rect 490158 687218 495522 687454
rect 495758 687218 501122 687454
rect 501358 687218 506722 687454
rect 506958 687218 510322 687454
rect 510558 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 85922 687134
rect 86158 686898 88522 687134
rect 88758 686898 95722 687134
rect 95958 686898 102922 687134
rect 103158 686898 110122 687134
rect 110358 686898 117322 687134
rect 117558 686898 119922 687134
rect 120158 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 241162 687134
rect 241398 686898 243762 687134
rect 243998 686898 250962 687134
rect 251198 686898 258162 687134
rect 258398 686898 265362 687134
rect 265598 686898 272562 687134
rect 272798 686898 275162 687134
rect 275398 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 486322 687134
rect 486558 686898 489922 687134
rect 490158 686898 495522 687134
rect 495758 686898 501122 687134
rect 501358 686898 506722 687134
rect 506958 686898 510322 687134
rect 510558 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 84922 669454
rect 85158 669218 92122 669454
rect 92358 669218 99322 669454
rect 99558 669218 106522 669454
rect 106758 669218 113722 669454
rect 113958 669218 120922 669454
rect 121158 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 240162 669454
rect 240398 669218 247362 669454
rect 247598 669218 254562 669454
rect 254798 669218 261762 669454
rect 261998 669218 268962 669454
rect 269198 669218 276162 669454
rect 276398 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487122 669454
rect 487358 669218 492722 669454
rect 492958 669218 498322 669454
rect 498558 669218 503922 669454
rect 504158 669218 509522 669454
rect 509758 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 84922 669134
rect 85158 668898 92122 669134
rect 92358 668898 99322 669134
rect 99558 668898 106522 669134
rect 106758 668898 113722 669134
rect 113958 668898 120922 669134
rect 121158 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 240162 669134
rect 240398 668898 247362 669134
rect 247598 668898 254562 669134
rect 254798 668898 261762 669134
rect 261998 668898 268962 669134
rect 269198 668898 276162 669134
rect 276398 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487122 669134
rect 487358 668898 492722 669134
rect 492958 668898 498322 669134
rect 498558 668898 503922 669134
rect 504158 668898 509522 669134
rect 509758 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 79542 615454
rect 79778 615218 110262 615454
rect 110498 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 239450 615454
rect 239686 615218 270170 615454
rect 270406 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 478998 615454
rect 479234 615218 509718 615454
rect 509954 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 79542 615134
rect 79778 614898 110262 615134
rect 110498 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 239450 615134
rect 239686 614898 270170 615134
rect 270406 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 478998 615134
rect 479234 614898 509718 615134
rect 509954 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 94902 597454
rect 95138 597218 125622 597454
rect 125858 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 254810 597454
rect 255046 597218 285530 597454
rect 285766 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 494358 597454
rect 494594 597218 525078 597454
rect 525314 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 94902 597134
rect 95138 596898 125622 597134
rect 125858 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 254810 597134
rect 255046 596898 285530 597134
rect 285766 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 494358 597134
rect 494594 596898 525078 597134
rect 525314 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 79542 579454
rect 79778 579218 110262 579454
rect 110498 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 239450 579454
rect 239686 579218 270170 579454
rect 270406 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 478998 579454
rect 479234 579218 509718 579454
rect 509954 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 79542 579134
rect 79778 578898 110262 579134
rect 110498 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 239450 579134
rect 239686 578898 270170 579134
rect 270406 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 478998 579134
rect 479234 578898 509718 579134
rect 509954 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 92426 562054
rect 92662 561818 92746 562054
rect 92982 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 92426 561734
rect 92662 561498 92746 561734
rect 92982 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 21008 399454
rect 21244 399218 155376 399454
rect 155612 399218 181008 399454
rect 181244 399218 315376 399454
rect 315612 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 21008 399134
rect 21244 398898 155376 399134
rect 155612 398898 181008 399134
rect 181244 398898 315376 399134
rect 315612 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 20328 381454
rect 20564 381218 156056 381454
rect 156292 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 180328 381454
rect 180564 381218 316056 381454
rect 316292 381218 359610 381454
rect 359846 381218 390330 381454
rect 390566 381218 421050 381454
rect 421286 381218 451770 381454
rect 452006 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 20328 381134
rect 20564 380898 156056 381134
rect 156292 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 180328 381134
rect 180564 380898 316056 381134
rect 316292 380898 359610 381134
rect 359846 380898 390330 381134
rect 390566 380898 421050 381134
rect 421286 380898 451770 381134
rect 452006 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 21008 363454
rect 21244 363218 155376 363454
rect 155612 363218 181008 363454
rect 181244 363218 315376 363454
rect 315612 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 344250 363454
rect 344486 363218 374970 363454
rect 375206 363218 405690 363454
rect 405926 363218 436410 363454
rect 436646 363218 467130 363454
rect 467366 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 21008 363134
rect 21244 362898 155376 363134
rect 155612 362898 181008 363134
rect 181244 362898 315376 363134
rect 315612 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 344250 363134
rect 344486 362898 374970 363134
rect 375206 362898 405690 363134
rect 405926 362898 436410 363134
rect 436646 362898 467130 363134
rect 467366 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 20328 345454
rect 20564 345218 156056 345454
rect 156292 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 180328 345454
rect 180564 345218 316056 345454
rect 316292 345218 359610 345454
rect 359846 345218 390330 345454
rect 390566 345218 421050 345454
rect 421286 345218 451770 345454
rect 452006 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 20328 345134
rect 20564 344898 156056 345134
rect 156292 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 180328 345134
rect 180564 344898 316056 345134
rect 316292 344898 359610 345134
rect 359846 344898 390330 345134
rect 390566 344898 421050 345134
rect 421286 344898 451770 345134
rect 452006 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 523130 331174
rect 523366 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 553850 331174
rect 554086 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 523130 330854
rect 523366 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 553850 330854
rect 554086 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 21008 327454
rect 21244 327218 155376 327454
rect 155612 327218 181008 327454
rect 181244 327218 315376 327454
rect 315612 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 344250 327454
rect 344486 327218 374970 327454
rect 375206 327218 405690 327454
rect 405926 327218 436410 327454
rect 436646 327218 467130 327454
rect 467366 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 507770 327454
rect 508006 327218 538490 327454
rect 538726 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 569210 327454
rect 569446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 21008 327134
rect 21244 326898 155376 327134
rect 155612 326898 181008 327134
rect 181244 326898 315376 327134
rect 315612 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 344250 327134
rect 344486 326898 374970 327134
rect 375206 326898 405690 327134
rect 405926 326898 436410 327134
rect 436646 326898 467130 327134
rect 467366 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 507770 327134
rect 508006 326898 538490 327134
rect 538726 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 569210 327134
rect 569446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 359610 309454
rect 359846 309218 390330 309454
rect 390566 309218 421050 309454
rect 421286 309218 451770 309454
rect 452006 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 359610 309134
rect 359846 308898 390330 309134
rect 390566 308898 421050 309134
rect 421286 308898 451770 309134
rect 452006 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect 30954 301674 283574 301706
rect 30954 301438 30986 301674
rect 31222 301438 31306 301674
rect 31542 301438 66986 301674
rect 67222 301438 67306 301674
rect 67542 301438 102986 301674
rect 103222 301438 103306 301674
rect 103542 301438 138986 301674
rect 139222 301438 139306 301674
rect 139542 301438 174986 301674
rect 175222 301438 175306 301674
rect 175542 301438 210986 301674
rect 211222 301438 211306 301674
rect 211542 301438 246986 301674
rect 247222 301438 247306 301674
rect 247542 301438 282986 301674
rect 283222 301438 283306 301674
rect 283542 301438 283574 301674
rect 30954 301354 283574 301438
rect 30954 301118 30986 301354
rect 31222 301118 31306 301354
rect 31542 301118 66986 301354
rect 67222 301118 67306 301354
rect 67542 301118 102986 301354
rect 103222 301118 103306 301354
rect 103542 301118 138986 301354
rect 139222 301118 139306 301354
rect 139542 301118 174986 301354
rect 175222 301118 175306 301354
rect 175542 301118 210986 301354
rect 211222 301118 211306 301354
rect 211542 301118 246986 301354
rect 247222 301118 247306 301354
rect 247542 301118 282986 301354
rect 283222 301118 283306 301354
rect 283542 301118 283574 301354
rect 30954 301086 283574 301118
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 31610 295174
rect 31846 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 62330 295174
rect 62566 294938 93050 295174
rect 93286 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 123770 295174
rect 124006 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 154490 295174
rect 154726 294938 185210 295174
rect 185446 294938 215930 295174
rect 216166 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 246650 295174
rect 246886 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 277370 295174
rect 277606 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 308090 295174
rect 308326 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 523130 295174
rect 523366 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 553850 295174
rect 554086 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 31610 294854
rect 31846 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 62330 294854
rect 62566 294618 93050 294854
rect 93286 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 123770 294854
rect 124006 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 154490 294854
rect 154726 294618 185210 294854
rect 185446 294618 215930 294854
rect 216166 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 246650 294854
rect 246886 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 277370 294854
rect 277606 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 308090 294854
rect 308326 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 523130 294854
rect 523366 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 553850 294854
rect 554086 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 16250 291454
rect 16486 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 46970 291454
rect 47206 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 139130 291454
rect 139366 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 169850 291454
rect 170086 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 200570 291454
rect 200806 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 231290 291454
rect 231526 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 262010 291454
rect 262246 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 344250 291454
rect 344486 291218 374970 291454
rect 375206 291218 405690 291454
rect 405926 291218 436410 291454
rect 436646 291218 467130 291454
rect 467366 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 507770 291454
rect 508006 291218 538490 291454
rect 538726 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 569210 291454
rect 569446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 16250 291134
rect 16486 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 46970 291134
rect 47206 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 139130 291134
rect 139366 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 169850 291134
rect 170086 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 200570 291134
rect 200806 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 231290 291134
rect 231526 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 262010 291134
rect 262246 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 344250 291134
rect 344486 290898 374970 291134
rect 375206 290898 405690 291134
rect 405926 290898 436410 291134
rect 436646 290898 467130 291134
rect 467366 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 507770 291134
rect 508006 290898 538490 291134
rect 538726 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 569210 291134
rect 569446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 20328 273454
rect 20564 273218 156056 273454
rect 156292 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 180328 273454
rect 180564 273218 316056 273454
rect 316292 273218 359610 273454
rect 359846 273218 390330 273454
rect 390566 273218 421050 273454
rect 421286 273218 451770 273454
rect 452006 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 20328 273134
rect 20564 272898 156056 273134
rect 156292 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 180328 273134
rect 180564 272898 316056 273134
rect 316292 272898 359610 273134
rect 359846 272898 390330 273134
rect 390566 272898 421050 273134
rect 421286 272898 451770 273134
rect 452006 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 523130 259174
rect 523366 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 553850 259174
rect 554086 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 523130 258854
rect 523366 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 553850 258854
rect 554086 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 21008 255454
rect 21244 255218 155376 255454
rect 155612 255218 181008 255454
rect 181244 255218 315376 255454
rect 315612 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 354170 255454
rect 354406 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 384890 255454
rect 385126 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 415610 255454
rect 415846 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 446330 255454
rect 446566 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 477050 255454
rect 477286 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 507770 255454
rect 508006 255218 538490 255454
rect 538726 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 569210 255454
rect 569446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 21008 255134
rect 21244 254898 155376 255134
rect 155612 254898 181008 255134
rect 181244 254898 315376 255134
rect 315612 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 354170 255134
rect 354406 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 384890 255134
rect 385126 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 415610 255134
rect 415846 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 446330 255134
rect 446566 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 477050 255134
rect 477286 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 507770 255134
rect 508006 254898 538490 255134
rect 538726 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 569210 255134
rect 569446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 20328 237454
rect 20564 237218 156056 237454
rect 156292 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 180328 237454
rect 180564 237218 316056 237454
rect 316292 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 20328 237134
rect 20564 236898 156056 237134
rect 156292 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 180328 237134
rect 180564 236898 316056 237134
rect 316292 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 338810 223174
rect 339046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 369530 223174
rect 369766 222938 400250 223174
rect 400486 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 430970 223174
rect 431206 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 461690 223174
rect 461926 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 492410 223174
rect 492646 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 523130 223174
rect 523366 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 553850 223174
rect 554086 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 338810 222854
rect 339046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 369530 222854
rect 369766 222618 400250 222854
rect 400486 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 430970 222854
rect 431206 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 461690 222854
rect 461926 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 492410 222854
rect 492646 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 523130 222854
rect 523366 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 553850 222854
rect 554086 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 21008 219454
rect 21244 219218 155376 219454
rect 155612 219218 181008 219454
rect 181244 219218 315376 219454
rect 315612 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 354170 219454
rect 354406 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 384890 219454
rect 385126 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 415610 219454
rect 415846 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 446330 219454
rect 446566 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 477050 219454
rect 477286 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 507770 219454
rect 508006 219218 538490 219454
rect 538726 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 569210 219454
rect 569446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 21008 219134
rect 21244 218898 155376 219134
rect 155612 218898 181008 219134
rect 181244 218898 315376 219134
rect 315612 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 354170 219134
rect 354406 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 384890 219134
rect 385126 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 415610 219134
rect 415846 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 446330 219134
rect 446566 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 477050 219134
rect 477286 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 507770 219134
rect 508006 218898 538490 219134
rect 538726 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 569210 219134
rect 569446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 31610 187174
rect 31846 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 62330 187174
rect 62566 186938 93050 187174
rect 93286 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 123770 187174
rect 124006 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 154490 187174
rect 154726 186938 185210 187174
rect 185446 186938 215930 187174
rect 216166 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 246650 187174
rect 246886 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 277370 187174
rect 277606 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 308090 187174
rect 308326 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 338810 187174
rect 339046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 369530 187174
rect 369766 186938 400250 187174
rect 400486 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 430970 187174
rect 431206 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 461690 187174
rect 461926 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 492410 187174
rect 492646 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 523130 187174
rect 523366 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 553850 187174
rect 554086 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 31610 186854
rect 31846 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 62330 186854
rect 62566 186618 93050 186854
rect 93286 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 123770 186854
rect 124006 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 154490 186854
rect 154726 186618 185210 186854
rect 185446 186618 215930 186854
rect 216166 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 246650 186854
rect 246886 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 277370 186854
rect 277606 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 308090 186854
rect 308326 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 338810 186854
rect 339046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 369530 186854
rect 369766 186618 400250 186854
rect 400486 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 430970 186854
rect 431206 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 461690 186854
rect 461926 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 492410 186854
rect 492646 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 523130 186854
rect 523366 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 553850 186854
rect 554086 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 16250 183454
rect 16486 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 46970 183454
rect 47206 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 139130 183454
rect 139366 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 169850 183454
rect 170086 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 200570 183454
rect 200806 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 231290 183454
rect 231526 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 262010 183454
rect 262246 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 354170 183454
rect 354406 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 384890 183454
rect 385126 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 415610 183454
rect 415846 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 446330 183454
rect 446566 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 477050 183454
rect 477286 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 507770 183454
rect 508006 183218 538490 183454
rect 538726 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 569210 183454
rect 569446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 16250 183134
rect 16486 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 46970 183134
rect 47206 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 139130 183134
rect 139366 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 169850 183134
rect 170086 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 200570 183134
rect 200806 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 231290 183134
rect 231526 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 262010 183134
rect 262246 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 354170 183134
rect 354406 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 384890 183134
rect 385126 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 415610 183134
rect 415846 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 446330 183134
rect 446566 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 477050 183134
rect 477286 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 507770 183134
rect 508006 182898 538490 183134
rect 538726 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 569210 183134
rect 569446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 31610 151174
rect 31846 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 62330 151174
rect 62566 150938 93050 151174
rect 93286 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 123770 151174
rect 124006 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 154490 151174
rect 154726 150938 185210 151174
rect 185446 150938 215930 151174
rect 216166 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 246650 151174
rect 246886 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 277370 151174
rect 277606 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 308090 151174
rect 308326 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 338810 151174
rect 339046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 369530 151174
rect 369766 150938 400250 151174
rect 400486 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 430970 151174
rect 431206 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 461690 151174
rect 461926 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 492410 151174
rect 492646 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 523130 151174
rect 523366 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 553850 151174
rect 554086 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 31610 150854
rect 31846 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 62330 150854
rect 62566 150618 93050 150854
rect 93286 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 123770 150854
rect 124006 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 154490 150854
rect 154726 150618 185210 150854
rect 185446 150618 215930 150854
rect 216166 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 246650 150854
rect 246886 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 277370 150854
rect 277606 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 308090 150854
rect 308326 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 338810 150854
rect 339046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 369530 150854
rect 369766 150618 400250 150854
rect 400486 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 430970 150854
rect 431206 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 461690 150854
rect 461926 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 492410 150854
rect 492646 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 523130 150854
rect 523366 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 553850 150854
rect 554086 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 16250 147454
rect 16486 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 46970 147454
rect 47206 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 139130 147454
rect 139366 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 169850 147454
rect 170086 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 200570 147454
rect 200806 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 231290 147454
rect 231526 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 262010 147454
rect 262246 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 354170 147454
rect 354406 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 384890 147454
rect 385126 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 415610 147454
rect 415846 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 446330 147454
rect 446566 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 477050 147454
rect 477286 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 507770 147454
rect 508006 147218 538490 147454
rect 538726 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 569210 147454
rect 569446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 16250 147134
rect 16486 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 46970 147134
rect 47206 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 139130 147134
rect 139366 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 169850 147134
rect 170086 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 200570 147134
rect 200806 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 231290 147134
rect 231526 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 262010 147134
rect 262246 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 354170 147134
rect 354406 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 384890 147134
rect 385126 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 415610 147134
rect 415846 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 446330 147134
rect 446566 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 477050 147134
rect 477286 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 507770 147134
rect 508006 146898 538490 147134
rect 538726 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 569210 147134
rect 569446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 31610 115174
rect 31846 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 62330 115174
rect 62566 114938 93050 115174
rect 93286 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 123770 115174
rect 124006 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 154490 115174
rect 154726 114938 185210 115174
rect 185446 114938 215930 115174
rect 216166 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 246650 115174
rect 246886 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 277370 115174
rect 277606 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 308090 115174
rect 308326 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 338810 115174
rect 339046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 369530 115174
rect 369766 114938 400250 115174
rect 400486 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 430970 115174
rect 431206 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 461690 115174
rect 461926 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 492410 115174
rect 492646 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 523130 115174
rect 523366 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 553850 115174
rect 554086 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 31610 114854
rect 31846 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 62330 114854
rect 62566 114618 93050 114854
rect 93286 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 123770 114854
rect 124006 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 154490 114854
rect 154726 114618 185210 114854
rect 185446 114618 215930 114854
rect 216166 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 246650 114854
rect 246886 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 277370 114854
rect 277606 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 308090 114854
rect 308326 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 338810 114854
rect 339046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 369530 114854
rect 369766 114618 400250 114854
rect 400486 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 430970 114854
rect 431206 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 461690 114854
rect 461926 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 492410 114854
rect 492646 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 523130 114854
rect 523366 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 553850 114854
rect 554086 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 16250 111454
rect 16486 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 46970 111454
rect 47206 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 139130 111454
rect 139366 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 169850 111454
rect 170086 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 200570 111454
rect 200806 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 231290 111454
rect 231526 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 262010 111454
rect 262246 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 354170 111454
rect 354406 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 384890 111454
rect 385126 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 415610 111454
rect 415846 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 446330 111454
rect 446566 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 477050 111454
rect 477286 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 507770 111454
rect 508006 111218 538490 111454
rect 538726 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 569210 111454
rect 569446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 16250 111134
rect 16486 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 46970 111134
rect 47206 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 139130 111134
rect 139366 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 169850 111134
rect 170086 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 200570 111134
rect 200806 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 231290 111134
rect 231526 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 262010 111134
rect 262246 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 354170 111134
rect 354406 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 384890 111134
rect 385126 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 415610 111134
rect 415846 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 446330 111134
rect 446566 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 477050 111134
rect 477286 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 507770 111134
rect 508006 110898 538490 111134
rect 538726 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 569210 111134
rect 569446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 31610 79174
rect 31846 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 62330 79174
rect 62566 78938 93050 79174
rect 93286 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 123770 79174
rect 124006 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 154490 79174
rect 154726 78938 185210 79174
rect 185446 78938 215930 79174
rect 216166 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 246650 79174
rect 246886 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 277370 79174
rect 277606 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 308090 79174
rect 308326 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 338810 79174
rect 339046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 369530 79174
rect 369766 78938 400250 79174
rect 400486 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 430970 79174
rect 431206 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 461690 79174
rect 461926 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 492410 79174
rect 492646 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 523130 79174
rect 523366 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 553850 79174
rect 554086 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 31610 78854
rect 31846 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 62330 78854
rect 62566 78618 93050 78854
rect 93286 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 123770 78854
rect 124006 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 154490 78854
rect 154726 78618 185210 78854
rect 185446 78618 215930 78854
rect 216166 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 246650 78854
rect 246886 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 277370 78854
rect 277606 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 308090 78854
rect 308326 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 338810 78854
rect 339046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 369530 78854
rect 369766 78618 400250 78854
rect 400486 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 430970 78854
rect 431206 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 461690 78854
rect 461926 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 492410 78854
rect 492646 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 523130 78854
rect 523366 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 553850 78854
rect 554086 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 16250 75454
rect 16486 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 46970 75454
rect 47206 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 139130 75454
rect 139366 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 169850 75454
rect 170086 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 200570 75454
rect 200806 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 231290 75454
rect 231526 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 262010 75454
rect 262246 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 354170 75454
rect 354406 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 384890 75454
rect 385126 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 415610 75454
rect 415846 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 446330 75454
rect 446566 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 477050 75454
rect 477286 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 507770 75454
rect 508006 75218 538490 75454
rect 538726 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 569210 75454
rect 569446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 16250 75134
rect 16486 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 46970 75134
rect 47206 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 139130 75134
rect 139366 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 169850 75134
rect 170086 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 200570 75134
rect 200806 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 231290 75134
rect 231526 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 262010 75134
rect 262246 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 354170 75134
rect 354406 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 384890 75134
rect 385126 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 415610 75134
rect 415846 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 446330 75134
rect 446566 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 477050 75134
rect 477286 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 507770 75134
rect 508006 74898 538490 75134
rect 538726 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 569210 75134
rect 569446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 31610 43174
rect 31846 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 62330 43174
rect 62566 42938 93050 43174
rect 93286 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 123770 43174
rect 124006 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 154490 43174
rect 154726 42938 185210 43174
rect 185446 42938 215930 43174
rect 216166 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 246650 43174
rect 246886 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 277370 43174
rect 277606 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 308090 43174
rect 308326 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 338810 43174
rect 339046 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 369530 43174
rect 369766 42938 400250 43174
rect 400486 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 430970 43174
rect 431206 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 461690 43174
rect 461926 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 492410 43174
rect 492646 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 523130 43174
rect 523366 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 553850 43174
rect 554086 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 31610 42854
rect 31846 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 62330 42854
rect 62566 42618 93050 42854
rect 93286 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 123770 42854
rect 124006 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 154490 42854
rect 154726 42618 185210 42854
rect 185446 42618 215930 42854
rect 216166 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 246650 42854
rect 246886 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 277370 42854
rect 277606 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 308090 42854
rect 308326 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 338810 42854
rect 339046 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 369530 42854
rect 369766 42618 400250 42854
rect 400486 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 430970 42854
rect 431206 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 461690 42854
rect 461926 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 492410 42854
rect 492646 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 523130 42854
rect 523366 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 553850 42854
rect 554086 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 16250 39454
rect 16486 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 46970 39454
rect 47206 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 139130 39454
rect 139366 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 169850 39454
rect 170086 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 200570 39454
rect 200806 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 231290 39454
rect 231526 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 262010 39454
rect 262246 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 354170 39454
rect 354406 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 384890 39454
rect 385126 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 415610 39454
rect 415846 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 446330 39454
rect 446566 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 477050 39454
rect 477286 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 507770 39454
rect 508006 39218 538490 39454
rect 538726 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 569210 39454
rect 569446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 16250 39134
rect 16486 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 46970 39134
rect 47206 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 139130 39134
rect 139366 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 169850 39134
rect 170086 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 200570 39134
rect 200806 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 231290 39134
rect 231526 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 262010 39134
rect 262246 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 354170 39134
rect 354406 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 384890 39134
rect 385126 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 415610 39134
rect 415846 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 446330 39134
rect 446566 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 477050 39134
rect 477286 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 507770 39134
rect 508006 38898 538490 39134
rect 538726 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 569210 39134
rect 569446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 31610 7174
rect 31846 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 62330 7174
rect 62566 6938 93050 7174
rect 93286 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 123770 7174
rect 124006 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 154490 7174
rect 154726 6938 185210 7174
rect 185446 6938 215930 7174
rect 216166 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 246650 7174
rect 246886 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 277370 7174
rect 277606 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 308090 7174
rect 308326 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 338810 7174
rect 339046 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 369530 7174
rect 369766 6938 400250 7174
rect 400486 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 430970 7174
rect 431206 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 461690 7174
rect 461926 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 492410 7174
rect 492646 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 523130 7174
rect 523366 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 553850 7174
rect 554086 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 31610 6854
rect 31846 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 62330 6854
rect 62566 6618 93050 6854
rect 93286 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 123770 6854
rect 124006 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 154490 6854
rect 154726 6618 185210 6854
rect 185446 6618 215930 6854
rect 216166 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 246650 6854
rect 246886 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 277370 6854
rect 277606 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 308090 6854
rect 308326 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 338810 6854
rect 339046 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 369530 6854
rect 369766 6618 400250 6854
rect 400486 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 430970 6854
rect 431206 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 461690 6854
rect 461926 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 492410 6854
rect 492646 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 523130 6854
rect 523366 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 553850 6854
rect 554086 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  mem_0
timestamp 1637984468
transform 1 0 20000 0 1 204000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  mem_1
timestamp 1637984468
transform 1 0 20000 0 1 322400
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  mem_2
timestamp 1637984468
transform 1 0 180000 0 1 204000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  mem_3
timestamp 1637984468
transform 1 0 180000 0 1 322400
box 0 0 136620 83308
use vco_adc_wrapper  vco_adc_wrapper_1
timestamp 1637984468
transform 1 0 340000 0 1 258000
box 0 0 140000 140000
use vco_adc  vco_adc_2
timestamp 1637984468
transform 1 0 75292 0 1 575820
box 0 0 53162 54000
use vco_adc  vco_adc_1
timestamp 1637984468
transform 1 0 235200 0 1 575820
box 0 0 53162 54000
use vco_adc  vco_adc_0
timestamp 1637984468
transform 1 0 474748 0 1 575820
box 0 0 53162 54000
use vco_r100  vco_2
timestamp 1637984468
transform 1 0 84840 0 1 667600
box 0 0 36702 21000
use vco  vco_1
timestamp 1637984468
transform 1 0 240080 0 1 667600
box 0 0 36602 21000
use vco_w6_r100  vco_0
timestamp 1637984468
transform 1 0 486240 0 1 667600
box 0 0 24610 21000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 202000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 256000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 256000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 256000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 256000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 289308 38414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 289308 74414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 289308 110414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 289308 146414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 289308 182414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 289308 218414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 289308 254414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 289308 290414 320400 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 407708 74414 573820 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 407708 110414 573820 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 407708 254414 573820 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 407708 290414 573820 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 573820 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 631820 110414 665600 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 631820 254414 665600 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 631820 506414 665600 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 407708 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 631820 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 690600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 407708 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 407708 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 407708 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 690600 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 631820 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 400000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 400000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 400000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 400000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 690600 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 202000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 256000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 256000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 256000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 256000 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 289308 42134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 289308 78134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 289308 114134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 289308 150134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 289308 186134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 289308 222134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 289308 258134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 289308 294134 320400 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 407708 78134 573820 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 407708 114134 573820 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 407708 258134 573820 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 400000 474134 573820 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 573820 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 631820 114134 665600 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 631820 258134 665600 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 631820 510134 665600 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 407708 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 631820 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 690600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 407708 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 407708 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 407708 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 690600 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 407708 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 400000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 400000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 400000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 631820 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 690600 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 202000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 256000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 256000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 256000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 256000 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 289308 45854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 289308 81854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 289308 117854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 289308 153854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 289308 189854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 289308 225854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 289308 261854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 289308 297854 320400 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 407708 81854 573820 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 407708 117854 573820 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 407708 261854 573820 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 400000 477854 573820 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 573820 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 631820 117854 665600 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 631820 261854 665600 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 407708 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 631820 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 690600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 407708 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 407708 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 407708 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 690600 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 407708 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 400000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 400000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 400000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 631820 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 631820 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 202000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 256000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 256000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 256000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 256000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 289308 49574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 289308 85574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 289308 121574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 289308 157574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 289308 193574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 289308 229574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 289308 265574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 289308 301574 320400 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 407708 85574 573820 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 407708 121574 573820 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 407708 265574 573820 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 400000 481574 573820 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 573820 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 631820 85574 665600 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 631820 121574 665600 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 631820 265574 665600 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 407708 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 690600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 690600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 407708 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 407708 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 407708 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 690600 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 407708 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 400000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 400000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 400000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 631820 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 631820 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 202000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 256000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 256000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 256000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 256000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 289308 27854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 289308 63854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 289308 99854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 289308 135854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 289308 207854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 289308 243854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 289308 279854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 289308 315854 320400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 407708 99854 573820 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 407708 243854 573820 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 407708 279854 573820 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 573820 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 631820 99854 665600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 631820 243854 665600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 631820 495854 665600 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 407708 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 407708 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 690600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 407708 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 407708 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 690600 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 631820 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 407708 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 400000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 400000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 400000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 400000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 690600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 30954 301086 283574 301706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 202000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 256000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 256000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 256000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 256000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 289308 31574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 289308 67574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 289308 103574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 289308 139574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 289308 211574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 289308 247574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 289308 283574 320400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 407708 103574 573820 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 407708 247574 573820 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 407708 283574 573820 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 573820 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 631820 103574 665600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 631820 247574 665600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 631820 499574 665600 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 407708 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 407708 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 690600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 407708 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 407708 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 690600 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 631820 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 400000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 400000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 400000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 400000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 690600 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 202000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 256000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 256000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 256000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 256000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 289308 20414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 289308 56414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 289308 92414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 289308 128414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 289308 200414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 289308 236414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 289308 272414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 289308 308414 320400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 407708 92414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 407708 128414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 407708 236414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 407708 272414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 573820 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 631820 92414 665600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 631820 272414 665600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 631820 488414 665600 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 407708 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 407708 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 690600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 631820 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 407708 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 631820 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 690600 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 407708 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 400000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 400000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 400000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 400000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 690600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 631820 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 202000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 256000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 256000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 256000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 256000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 289308 24134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 289308 60134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 289308 96134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 289308 132134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 289308 204134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 289308 240134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 289308 276134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 289308 312134 320400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 407708 96134 573820 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 407708 240134 573820 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 407708 276134 573820 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 573820 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 573820 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 631820 96134 665600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 631820 240134 665600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 631820 276134 665600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 631820 492134 665600 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 407708 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 407708 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 690600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 407708 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 407708 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 690600 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 690600 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 407708 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 400000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 400000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 400000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 400000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 690600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 631820 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
