magic
tech sky130A
magscale 1 2
timestamp 1695114543
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 934 1776 139090 137680
<< metal2 >>
rect 3146 139200 3202 140000
rect 4158 139200 4214 140000
rect 5170 139200 5226 140000
rect 6182 139200 6238 140000
rect 7194 139200 7250 140000
rect 8206 139200 8262 140000
rect 9218 139200 9274 140000
rect 10230 139200 10286 140000
rect 11242 139200 11298 140000
rect 12254 139200 12310 140000
rect 13266 139200 13322 140000
rect 14278 139200 14334 140000
rect 15290 139200 15346 140000
rect 16302 139200 16358 140000
rect 17314 139200 17370 140000
rect 18326 139200 18382 140000
rect 19338 139200 19394 140000
rect 20350 139200 20406 140000
rect 21362 139200 21418 140000
rect 22374 139200 22430 140000
rect 23386 139200 23442 140000
rect 24398 139200 24454 140000
rect 25410 139200 25466 140000
rect 26422 139200 26478 140000
rect 27434 139200 27490 140000
rect 28446 139200 28502 140000
rect 29458 139200 29514 140000
rect 30470 139200 30526 140000
rect 31482 139200 31538 140000
rect 32494 139200 32550 140000
rect 33506 139200 33562 140000
rect 34518 139200 34574 140000
rect 35530 139200 35586 140000
rect 36542 139200 36598 140000
rect 37554 139200 37610 140000
rect 38566 139200 38622 140000
rect 39578 139200 39634 140000
rect 40590 139200 40646 140000
rect 41602 139200 41658 140000
rect 42614 139200 42670 140000
rect 43626 139200 43682 140000
rect 44638 139200 44694 140000
rect 45650 139200 45706 140000
rect 46662 139200 46718 140000
rect 47674 139200 47730 140000
rect 48686 139200 48742 140000
rect 49698 139200 49754 140000
rect 50710 139200 50766 140000
rect 51722 139200 51778 140000
rect 52734 139200 52790 140000
rect 53746 139200 53802 140000
rect 54758 139200 54814 140000
rect 55770 139200 55826 140000
rect 56782 139200 56838 140000
rect 57794 139200 57850 140000
rect 58806 139200 58862 140000
rect 59818 139200 59874 140000
rect 60830 139200 60886 140000
rect 61842 139200 61898 140000
rect 62854 139200 62910 140000
rect 63866 139200 63922 140000
rect 64878 139200 64934 140000
rect 65890 139200 65946 140000
rect 66902 139200 66958 140000
rect 67914 139200 67970 140000
rect 68926 139200 68982 140000
rect 69938 139200 69994 140000
rect 70950 139200 71006 140000
rect 71962 139200 72018 140000
rect 72974 139200 73030 140000
rect 73986 139200 74042 140000
rect 74998 139200 75054 140000
rect 76010 139200 76066 140000
rect 77022 139200 77078 140000
rect 78034 139200 78090 140000
rect 79046 139200 79102 140000
rect 80058 139200 80114 140000
rect 81070 139200 81126 140000
rect 82082 139200 82138 140000
rect 83094 139200 83150 140000
rect 84106 139200 84162 140000
rect 85118 139200 85174 140000
rect 86130 139200 86186 140000
rect 87142 139200 87198 140000
rect 88154 139200 88210 140000
rect 89166 139200 89222 140000
rect 90178 139200 90234 140000
rect 91190 139200 91246 140000
rect 92202 139200 92258 140000
rect 93214 139200 93270 140000
rect 94226 139200 94282 140000
rect 95238 139200 95294 140000
rect 96250 139200 96306 140000
rect 97262 139200 97318 140000
rect 98274 139200 98330 140000
rect 99286 139200 99342 140000
rect 100298 139200 100354 140000
rect 101310 139200 101366 140000
rect 102322 139200 102378 140000
rect 103334 139200 103390 140000
rect 104346 139200 104402 140000
rect 105358 139200 105414 140000
rect 106370 139200 106426 140000
rect 107382 139200 107438 140000
rect 108394 139200 108450 140000
rect 109406 139200 109462 140000
rect 110418 139200 110474 140000
rect 111430 139200 111486 140000
rect 112442 139200 112498 140000
rect 113454 139200 113510 140000
rect 114466 139200 114522 140000
rect 115478 139200 115534 140000
rect 116490 139200 116546 140000
rect 117502 139200 117558 140000
rect 118514 139200 118570 140000
rect 119526 139200 119582 140000
rect 120538 139200 120594 140000
rect 121550 139200 121606 140000
rect 122562 139200 122618 140000
rect 123574 139200 123630 140000
rect 124586 139200 124642 140000
rect 125598 139200 125654 140000
rect 126610 139200 126666 140000
rect 127622 139200 127678 140000
rect 128634 139200 128690 140000
rect 129646 139200 129702 140000
rect 130658 139200 130714 140000
rect 131670 139200 131726 140000
rect 132682 139200 132738 140000
rect 133694 139200 133750 140000
rect 134706 139200 134762 140000
rect 135718 139200 135774 140000
rect 136730 139200 136786 140000
rect 2318 0 2374 800
rect 3606 0 3662 800
rect 4894 0 4950 800
rect 6182 0 6238 800
rect 7470 0 7526 800
rect 8758 0 8814 800
rect 10046 0 10102 800
rect 11334 0 11390 800
rect 12622 0 12678 800
rect 13910 0 13966 800
rect 15198 0 15254 800
rect 16486 0 16542 800
rect 17774 0 17830 800
rect 19062 0 19118 800
rect 20350 0 20406 800
rect 21638 0 21694 800
rect 22926 0 22982 800
rect 24214 0 24270 800
rect 25502 0 25558 800
rect 26790 0 26846 800
rect 28078 0 28134 800
rect 29366 0 29422 800
rect 30654 0 30710 800
rect 31942 0 31998 800
rect 33230 0 33286 800
rect 34518 0 34574 800
rect 35806 0 35862 800
rect 37094 0 37150 800
rect 38382 0 38438 800
rect 39670 0 39726 800
rect 40958 0 41014 800
rect 42246 0 42302 800
rect 43534 0 43590 800
rect 44822 0 44878 800
rect 46110 0 46166 800
rect 47398 0 47454 800
rect 48686 0 48742 800
rect 49974 0 50030 800
rect 51262 0 51318 800
rect 52550 0 52606 800
rect 53838 0 53894 800
rect 55126 0 55182 800
rect 56414 0 56470 800
rect 57702 0 57758 800
rect 58990 0 59046 800
rect 60278 0 60334 800
rect 61566 0 61622 800
rect 62854 0 62910 800
rect 64142 0 64198 800
rect 65430 0 65486 800
rect 66718 0 66774 800
rect 68006 0 68062 800
rect 69294 0 69350 800
rect 70582 0 70638 800
rect 71870 0 71926 800
rect 73158 0 73214 800
rect 74446 0 74502 800
rect 75734 0 75790 800
rect 77022 0 77078 800
rect 78310 0 78366 800
rect 79598 0 79654 800
rect 80886 0 80942 800
rect 82174 0 82230 800
rect 83462 0 83518 800
rect 84750 0 84806 800
rect 86038 0 86094 800
rect 87326 0 87382 800
rect 88614 0 88670 800
rect 89902 0 89958 800
rect 91190 0 91246 800
rect 92478 0 92534 800
rect 93766 0 93822 800
rect 95054 0 95110 800
rect 96342 0 96398 800
rect 97630 0 97686 800
rect 98918 0 98974 800
rect 100206 0 100262 800
rect 101494 0 101550 800
rect 102782 0 102838 800
rect 104070 0 104126 800
rect 105358 0 105414 800
rect 106646 0 106702 800
rect 107934 0 107990 800
rect 109222 0 109278 800
rect 110510 0 110566 800
rect 111798 0 111854 800
rect 113086 0 113142 800
rect 114374 0 114430 800
rect 115662 0 115718 800
rect 116950 0 117006 800
rect 118238 0 118294 800
rect 119526 0 119582 800
rect 120814 0 120870 800
rect 122102 0 122158 800
rect 123390 0 123446 800
rect 124678 0 124734 800
rect 125966 0 126022 800
rect 127254 0 127310 800
rect 128542 0 128598 800
rect 129830 0 129886 800
rect 131118 0 131174 800
rect 132406 0 132462 800
rect 133694 0 133750 800
rect 134982 0 135038 800
rect 136270 0 136326 800
rect 137558 0 137614 800
<< obsm2 >>
rect 938 139144 3090 139346
rect 3258 139144 4102 139346
rect 4270 139144 5114 139346
rect 5282 139144 6126 139346
rect 6294 139144 7138 139346
rect 7306 139144 8150 139346
rect 8318 139144 9162 139346
rect 9330 139144 10174 139346
rect 10342 139144 11186 139346
rect 11354 139144 12198 139346
rect 12366 139144 13210 139346
rect 13378 139144 14222 139346
rect 14390 139144 15234 139346
rect 15402 139144 16246 139346
rect 16414 139144 17258 139346
rect 17426 139144 18270 139346
rect 18438 139144 19282 139346
rect 19450 139144 20294 139346
rect 20462 139144 21306 139346
rect 21474 139144 22318 139346
rect 22486 139144 23330 139346
rect 23498 139144 24342 139346
rect 24510 139144 25354 139346
rect 25522 139144 26366 139346
rect 26534 139144 27378 139346
rect 27546 139144 28390 139346
rect 28558 139144 29402 139346
rect 29570 139144 30414 139346
rect 30582 139144 31426 139346
rect 31594 139144 32438 139346
rect 32606 139144 33450 139346
rect 33618 139144 34462 139346
rect 34630 139144 35474 139346
rect 35642 139144 36486 139346
rect 36654 139144 37498 139346
rect 37666 139144 38510 139346
rect 38678 139144 39522 139346
rect 39690 139144 40534 139346
rect 40702 139144 41546 139346
rect 41714 139144 42558 139346
rect 42726 139144 43570 139346
rect 43738 139144 44582 139346
rect 44750 139144 45594 139346
rect 45762 139144 46606 139346
rect 46774 139144 47618 139346
rect 47786 139144 48630 139346
rect 48798 139144 49642 139346
rect 49810 139144 50654 139346
rect 50822 139144 51666 139346
rect 51834 139144 52678 139346
rect 52846 139144 53690 139346
rect 53858 139144 54702 139346
rect 54870 139144 55714 139346
rect 55882 139144 56726 139346
rect 56894 139144 57738 139346
rect 57906 139144 58750 139346
rect 58918 139144 59762 139346
rect 59930 139144 60774 139346
rect 60942 139144 61786 139346
rect 61954 139144 62798 139346
rect 62966 139144 63810 139346
rect 63978 139144 64822 139346
rect 64990 139144 65834 139346
rect 66002 139144 66846 139346
rect 67014 139144 67858 139346
rect 68026 139144 68870 139346
rect 69038 139144 69882 139346
rect 70050 139144 70894 139346
rect 71062 139144 71906 139346
rect 72074 139144 72918 139346
rect 73086 139144 73930 139346
rect 74098 139144 74942 139346
rect 75110 139144 75954 139346
rect 76122 139144 76966 139346
rect 77134 139144 77978 139346
rect 78146 139144 78990 139346
rect 79158 139144 80002 139346
rect 80170 139144 81014 139346
rect 81182 139144 82026 139346
rect 82194 139144 83038 139346
rect 83206 139144 84050 139346
rect 84218 139144 85062 139346
rect 85230 139144 86074 139346
rect 86242 139144 87086 139346
rect 87254 139144 88098 139346
rect 88266 139144 89110 139346
rect 89278 139144 90122 139346
rect 90290 139144 91134 139346
rect 91302 139144 92146 139346
rect 92314 139144 93158 139346
rect 93326 139144 94170 139346
rect 94338 139144 95182 139346
rect 95350 139144 96194 139346
rect 96362 139144 97206 139346
rect 97374 139144 98218 139346
rect 98386 139144 99230 139346
rect 99398 139144 100242 139346
rect 100410 139144 101254 139346
rect 101422 139144 102266 139346
rect 102434 139144 103278 139346
rect 103446 139144 104290 139346
rect 104458 139144 105302 139346
rect 105470 139144 106314 139346
rect 106482 139144 107326 139346
rect 107494 139144 108338 139346
rect 108506 139144 109350 139346
rect 109518 139144 110362 139346
rect 110530 139144 111374 139346
rect 111542 139144 112386 139346
rect 112554 139144 113398 139346
rect 113566 139144 114410 139346
rect 114578 139144 115422 139346
rect 115590 139144 116434 139346
rect 116602 139144 117446 139346
rect 117614 139144 118458 139346
rect 118626 139144 119470 139346
rect 119638 139144 120482 139346
rect 120650 139144 121494 139346
rect 121662 139144 122506 139346
rect 122674 139144 123518 139346
rect 123686 139144 124530 139346
rect 124698 139144 125542 139346
rect 125710 139144 126554 139346
rect 126722 139144 127566 139346
rect 127734 139144 128578 139346
rect 128746 139144 129590 139346
rect 129758 139144 130602 139346
rect 130770 139144 131614 139346
rect 131782 139144 132626 139346
rect 132794 139144 133638 139346
rect 133806 139144 134650 139346
rect 134818 139144 135662 139346
rect 135830 139144 136674 139346
rect 136842 139144 139086 139346
rect 938 856 139086 139144
rect 938 734 2262 856
rect 2430 734 3550 856
rect 3718 734 4838 856
rect 5006 734 6126 856
rect 6294 734 7414 856
rect 7582 734 8702 856
rect 8870 734 9990 856
rect 10158 734 11278 856
rect 11446 734 12566 856
rect 12734 734 13854 856
rect 14022 734 15142 856
rect 15310 734 16430 856
rect 16598 734 17718 856
rect 17886 734 19006 856
rect 19174 734 20294 856
rect 20462 734 21582 856
rect 21750 734 22870 856
rect 23038 734 24158 856
rect 24326 734 25446 856
rect 25614 734 26734 856
rect 26902 734 28022 856
rect 28190 734 29310 856
rect 29478 734 30598 856
rect 30766 734 31886 856
rect 32054 734 33174 856
rect 33342 734 34462 856
rect 34630 734 35750 856
rect 35918 734 37038 856
rect 37206 734 38326 856
rect 38494 734 39614 856
rect 39782 734 40902 856
rect 41070 734 42190 856
rect 42358 734 43478 856
rect 43646 734 44766 856
rect 44934 734 46054 856
rect 46222 734 47342 856
rect 47510 734 48630 856
rect 48798 734 49918 856
rect 50086 734 51206 856
rect 51374 734 52494 856
rect 52662 734 53782 856
rect 53950 734 55070 856
rect 55238 734 56358 856
rect 56526 734 57646 856
rect 57814 734 58934 856
rect 59102 734 60222 856
rect 60390 734 61510 856
rect 61678 734 62798 856
rect 62966 734 64086 856
rect 64254 734 65374 856
rect 65542 734 66662 856
rect 66830 734 67950 856
rect 68118 734 69238 856
rect 69406 734 70526 856
rect 70694 734 71814 856
rect 71982 734 73102 856
rect 73270 734 74390 856
rect 74558 734 75678 856
rect 75846 734 76966 856
rect 77134 734 78254 856
rect 78422 734 79542 856
rect 79710 734 80830 856
rect 80998 734 82118 856
rect 82286 734 83406 856
rect 83574 734 84694 856
rect 84862 734 85982 856
rect 86150 734 87270 856
rect 87438 734 88558 856
rect 88726 734 89846 856
rect 90014 734 91134 856
rect 91302 734 92422 856
rect 92590 734 93710 856
rect 93878 734 94998 856
rect 95166 734 96286 856
rect 96454 734 97574 856
rect 97742 734 98862 856
rect 99030 734 100150 856
rect 100318 734 101438 856
rect 101606 734 102726 856
rect 102894 734 104014 856
rect 104182 734 105302 856
rect 105470 734 106590 856
rect 106758 734 107878 856
rect 108046 734 109166 856
rect 109334 734 110454 856
rect 110622 734 111742 856
rect 111910 734 113030 856
rect 113198 734 114318 856
rect 114486 734 115606 856
rect 115774 734 116894 856
rect 117062 734 118182 856
rect 118350 734 119470 856
rect 119638 734 120758 856
rect 120926 734 122046 856
rect 122214 734 123334 856
rect 123502 734 124622 856
rect 124790 734 125910 856
rect 126078 734 127198 856
rect 127366 734 128486 856
rect 128654 734 129774 856
rect 129942 734 131062 856
rect 131230 734 132350 856
rect 132518 734 133638 856
rect 133806 734 134926 856
rect 135094 734 136214 856
rect 136382 734 137502 856
rect 137670 734 139086 856
<< metal3 >>
rect 139200 136824 140000 136944
rect 139200 132200 140000 132320
rect 0 128936 800 129056
rect 0 128392 800 128512
rect 0 127848 800 127968
rect 139200 127576 140000 127696
rect 0 127304 800 127424
rect 0 126760 800 126880
rect 0 126216 800 126336
rect 0 125672 800 125792
rect 0 125128 800 125248
rect 0 124584 800 124704
rect 0 124040 800 124160
rect 0 123496 800 123616
rect 0 122952 800 123072
rect 139200 122952 140000 123072
rect 0 122408 800 122528
rect 0 121864 800 121984
rect 0 121320 800 121440
rect 0 120776 800 120896
rect 0 120232 800 120352
rect 0 119688 800 119808
rect 0 119144 800 119264
rect 0 118600 800 118720
rect 139200 118328 140000 118448
rect 0 118056 800 118176
rect 0 117512 800 117632
rect 0 116968 800 117088
rect 0 116424 800 116544
rect 0 115880 800 116000
rect 0 115336 800 115456
rect 0 114792 800 114912
rect 0 114248 800 114368
rect 0 113704 800 113824
rect 139200 113704 140000 113824
rect 0 113160 800 113280
rect 0 112616 800 112736
rect 0 112072 800 112192
rect 0 111528 800 111648
rect 0 110984 800 111104
rect 0 110440 800 110560
rect 0 109896 800 110016
rect 0 109352 800 109472
rect 139200 109080 140000 109200
rect 0 108808 800 108928
rect 0 108264 800 108384
rect 0 107720 800 107840
rect 0 107176 800 107296
rect 0 106632 800 106752
rect 0 106088 800 106208
rect 0 105544 800 105664
rect 0 105000 800 105120
rect 0 104456 800 104576
rect 139200 104456 140000 104576
rect 0 103912 800 104032
rect 0 103368 800 103488
rect 0 102824 800 102944
rect 0 102280 800 102400
rect 0 101736 800 101856
rect 0 101192 800 101312
rect 0 100648 800 100768
rect 0 100104 800 100224
rect 139200 99832 140000 99952
rect 0 99560 800 99680
rect 0 99016 800 99136
rect 0 98472 800 98592
rect 0 97928 800 98048
rect 0 97384 800 97504
rect 0 96840 800 96960
rect 0 96296 800 96416
rect 0 95752 800 95872
rect 0 95208 800 95328
rect 139200 95208 140000 95328
rect 0 94664 800 94784
rect 0 94120 800 94240
rect 0 93576 800 93696
rect 0 93032 800 93152
rect 0 92488 800 92608
rect 0 91944 800 92064
rect 0 91400 800 91520
rect 0 90856 800 90976
rect 139200 90584 140000 90704
rect 0 90312 800 90432
rect 0 89768 800 89888
rect 0 89224 800 89344
rect 0 88680 800 88800
rect 0 88136 800 88256
rect 0 87592 800 87712
rect 0 87048 800 87168
rect 0 86504 800 86624
rect 0 85960 800 86080
rect 139200 85960 140000 86080
rect 0 85416 800 85536
rect 0 84872 800 84992
rect 0 84328 800 84448
rect 0 83784 800 83904
rect 0 83240 800 83360
rect 0 82696 800 82816
rect 0 82152 800 82272
rect 0 81608 800 81728
rect 139200 81336 140000 81456
rect 0 81064 800 81184
rect 0 80520 800 80640
rect 0 79976 800 80096
rect 0 79432 800 79552
rect 0 78888 800 79008
rect 0 78344 800 78464
rect 0 77800 800 77920
rect 0 77256 800 77376
rect 0 76712 800 76832
rect 139200 76712 140000 76832
rect 0 76168 800 76288
rect 0 75624 800 75744
rect 0 75080 800 75200
rect 0 74536 800 74656
rect 0 73992 800 74112
rect 0 73448 800 73568
rect 0 72904 800 73024
rect 0 72360 800 72480
rect 139200 72088 140000 72208
rect 0 71816 800 71936
rect 0 71272 800 71392
rect 0 70728 800 70848
rect 0 70184 800 70304
rect 0 69640 800 69760
rect 0 69096 800 69216
rect 0 68552 800 68672
rect 0 68008 800 68128
rect 0 67464 800 67584
rect 139200 67464 140000 67584
rect 0 66920 800 67040
rect 0 66376 800 66496
rect 0 65832 800 65952
rect 0 65288 800 65408
rect 0 64744 800 64864
rect 0 64200 800 64320
rect 0 63656 800 63776
rect 0 63112 800 63232
rect 139200 62840 140000 62960
rect 0 62568 800 62688
rect 0 62024 800 62144
rect 0 61480 800 61600
rect 0 60936 800 61056
rect 0 60392 800 60512
rect 0 59848 800 59968
rect 0 59304 800 59424
rect 0 58760 800 58880
rect 0 58216 800 58336
rect 139200 58216 140000 58336
rect 0 57672 800 57792
rect 0 57128 800 57248
rect 0 56584 800 56704
rect 0 56040 800 56160
rect 0 55496 800 55616
rect 0 54952 800 55072
rect 0 54408 800 54528
rect 0 53864 800 53984
rect 139200 53592 140000 53712
rect 0 53320 800 53440
rect 0 52776 800 52896
rect 0 52232 800 52352
rect 0 51688 800 51808
rect 0 51144 800 51264
rect 0 50600 800 50720
rect 0 50056 800 50176
rect 0 49512 800 49632
rect 0 48968 800 49088
rect 139200 48968 140000 49088
rect 0 48424 800 48544
rect 0 47880 800 48000
rect 0 47336 800 47456
rect 0 46792 800 46912
rect 0 46248 800 46368
rect 0 45704 800 45824
rect 0 45160 800 45280
rect 0 44616 800 44736
rect 139200 44344 140000 44464
rect 0 44072 800 44192
rect 0 43528 800 43648
rect 0 42984 800 43104
rect 0 42440 800 42560
rect 0 41896 800 42016
rect 0 41352 800 41472
rect 0 40808 800 40928
rect 0 40264 800 40384
rect 0 39720 800 39840
rect 139200 39720 140000 39840
rect 0 39176 800 39296
rect 0 38632 800 38752
rect 0 38088 800 38208
rect 0 37544 800 37664
rect 0 37000 800 37120
rect 0 36456 800 36576
rect 0 35912 800 36032
rect 0 35368 800 35488
rect 139200 35096 140000 35216
rect 0 34824 800 34944
rect 0 34280 800 34400
rect 0 33736 800 33856
rect 0 33192 800 33312
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 0 31560 800 31680
rect 0 31016 800 31136
rect 0 30472 800 30592
rect 139200 30472 140000 30592
rect 0 29928 800 30048
rect 0 29384 800 29504
rect 0 28840 800 28960
rect 0 28296 800 28416
rect 0 27752 800 27872
rect 0 27208 800 27328
rect 0 26664 800 26784
rect 0 26120 800 26240
rect 139200 25848 140000 25968
rect 0 25576 800 25696
rect 0 25032 800 25152
rect 0 24488 800 24608
rect 0 23944 800 24064
rect 0 23400 800 23520
rect 0 22856 800 22976
rect 0 22312 800 22432
rect 0 21768 800 21888
rect 0 21224 800 21344
rect 139200 21224 140000 21344
rect 0 20680 800 20800
rect 0 20136 800 20256
rect 0 19592 800 19712
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 139200 16600 140000 16720
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 0 13608 800 13728
rect 0 13064 800 13184
rect 0 12520 800 12640
rect 0 11976 800 12096
rect 139200 11976 140000 12096
rect 0 11432 800 11552
rect 0 10888 800 11008
rect 139200 7352 140000 7472
rect 139200 2728 140000 2848
<< obsm3 >>
rect 798 137024 139200 137665
rect 798 136744 139120 137024
rect 798 132400 139200 136744
rect 798 132120 139120 132400
rect 798 129136 139200 132120
rect 880 128856 139200 129136
rect 798 128592 139200 128856
rect 880 128312 139200 128592
rect 798 128048 139200 128312
rect 880 127776 139200 128048
rect 880 127768 139120 127776
rect 798 127504 139120 127768
rect 880 127496 139120 127504
rect 880 127224 139200 127496
rect 798 126960 139200 127224
rect 880 126680 139200 126960
rect 798 126416 139200 126680
rect 880 126136 139200 126416
rect 798 125872 139200 126136
rect 880 125592 139200 125872
rect 798 125328 139200 125592
rect 880 125048 139200 125328
rect 798 124784 139200 125048
rect 880 124504 139200 124784
rect 798 124240 139200 124504
rect 880 123960 139200 124240
rect 798 123696 139200 123960
rect 880 123416 139200 123696
rect 798 123152 139200 123416
rect 880 122872 139120 123152
rect 798 122608 139200 122872
rect 880 122328 139200 122608
rect 798 122064 139200 122328
rect 880 121784 139200 122064
rect 798 121520 139200 121784
rect 880 121240 139200 121520
rect 798 120976 139200 121240
rect 880 120696 139200 120976
rect 798 120432 139200 120696
rect 880 120152 139200 120432
rect 798 119888 139200 120152
rect 880 119608 139200 119888
rect 798 119344 139200 119608
rect 880 119064 139200 119344
rect 798 118800 139200 119064
rect 880 118528 139200 118800
rect 880 118520 139120 118528
rect 798 118256 139120 118520
rect 880 118248 139120 118256
rect 880 117976 139200 118248
rect 798 117712 139200 117976
rect 880 117432 139200 117712
rect 798 117168 139200 117432
rect 880 116888 139200 117168
rect 798 116624 139200 116888
rect 880 116344 139200 116624
rect 798 116080 139200 116344
rect 880 115800 139200 116080
rect 798 115536 139200 115800
rect 880 115256 139200 115536
rect 798 114992 139200 115256
rect 880 114712 139200 114992
rect 798 114448 139200 114712
rect 880 114168 139200 114448
rect 798 113904 139200 114168
rect 880 113624 139120 113904
rect 798 113360 139200 113624
rect 880 113080 139200 113360
rect 798 112816 139200 113080
rect 880 112536 139200 112816
rect 798 112272 139200 112536
rect 880 111992 139200 112272
rect 798 111728 139200 111992
rect 880 111448 139200 111728
rect 798 111184 139200 111448
rect 880 110904 139200 111184
rect 798 110640 139200 110904
rect 880 110360 139200 110640
rect 798 110096 139200 110360
rect 880 109816 139200 110096
rect 798 109552 139200 109816
rect 880 109280 139200 109552
rect 880 109272 139120 109280
rect 798 109008 139120 109272
rect 880 109000 139120 109008
rect 880 108728 139200 109000
rect 798 108464 139200 108728
rect 880 108184 139200 108464
rect 798 107920 139200 108184
rect 880 107640 139200 107920
rect 798 107376 139200 107640
rect 880 107096 139200 107376
rect 798 106832 139200 107096
rect 880 106552 139200 106832
rect 798 106288 139200 106552
rect 880 106008 139200 106288
rect 798 105744 139200 106008
rect 880 105464 139200 105744
rect 798 105200 139200 105464
rect 880 104920 139200 105200
rect 798 104656 139200 104920
rect 880 104376 139120 104656
rect 798 104112 139200 104376
rect 880 103832 139200 104112
rect 798 103568 139200 103832
rect 880 103288 139200 103568
rect 798 103024 139200 103288
rect 880 102744 139200 103024
rect 798 102480 139200 102744
rect 880 102200 139200 102480
rect 798 101936 139200 102200
rect 880 101656 139200 101936
rect 798 101392 139200 101656
rect 880 101112 139200 101392
rect 798 100848 139200 101112
rect 880 100568 139200 100848
rect 798 100304 139200 100568
rect 880 100032 139200 100304
rect 880 100024 139120 100032
rect 798 99760 139120 100024
rect 880 99752 139120 99760
rect 880 99480 139200 99752
rect 798 99216 139200 99480
rect 880 98936 139200 99216
rect 798 98672 139200 98936
rect 880 98392 139200 98672
rect 798 98128 139200 98392
rect 880 97848 139200 98128
rect 798 97584 139200 97848
rect 880 97304 139200 97584
rect 798 97040 139200 97304
rect 880 96760 139200 97040
rect 798 96496 139200 96760
rect 880 96216 139200 96496
rect 798 95952 139200 96216
rect 880 95672 139200 95952
rect 798 95408 139200 95672
rect 880 95128 139120 95408
rect 798 94864 139200 95128
rect 880 94584 139200 94864
rect 798 94320 139200 94584
rect 880 94040 139200 94320
rect 798 93776 139200 94040
rect 880 93496 139200 93776
rect 798 93232 139200 93496
rect 880 92952 139200 93232
rect 798 92688 139200 92952
rect 880 92408 139200 92688
rect 798 92144 139200 92408
rect 880 91864 139200 92144
rect 798 91600 139200 91864
rect 880 91320 139200 91600
rect 798 91056 139200 91320
rect 880 90784 139200 91056
rect 880 90776 139120 90784
rect 798 90512 139120 90776
rect 880 90504 139120 90512
rect 880 90232 139200 90504
rect 798 89968 139200 90232
rect 880 89688 139200 89968
rect 798 89424 139200 89688
rect 880 89144 139200 89424
rect 798 88880 139200 89144
rect 880 88600 139200 88880
rect 798 88336 139200 88600
rect 880 88056 139200 88336
rect 798 87792 139200 88056
rect 880 87512 139200 87792
rect 798 87248 139200 87512
rect 880 86968 139200 87248
rect 798 86704 139200 86968
rect 880 86424 139200 86704
rect 798 86160 139200 86424
rect 880 85880 139120 86160
rect 798 85616 139200 85880
rect 880 85336 139200 85616
rect 798 85072 139200 85336
rect 880 84792 139200 85072
rect 798 84528 139200 84792
rect 880 84248 139200 84528
rect 798 83984 139200 84248
rect 880 83704 139200 83984
rect 798 83440 139200 83704
rect 880 83160 139200 83440
rect 798 82896 139200 83160
rect 880 82616 139200 82896
rect 798 82352 139200 82616
rect 880 82072 139200 82352
rect 798 81808 139200 82072
rect 880 81536 139200 81808
rect 880 81528 139120 81536
rect 798 81264 139120 81528
rect 880 81256 139120 81264
rect 880 80984 139200 81256
rect 798 80720 139200 80984
rect 880 80440 139200 80720
rect 798 80176 139200 80440
rect 880 79896 139200 80176
rect 798 79632 139200 79896
rect 880 79352 139200 79632
rect 798 79088 139200 79352
rect 880 78808 139200 79088
rect 798 78544 139200 78808
rect 880 78264 139200 78544
rect 798 78000 139200 78264
rect 880 77720 139200 78000
rect 798 77456 139200 77720
rect 880 77176 139200 77456
rect 798 76912 139200 77176
rect 880 76632 139120 76912
rect 798 76368 139200 76632
rect 880 76088 139200 76368
rect 798 75824 139200 76088
rect 880 75544 139200 75824
rect 798 75280 139200 75544
rect 880 75000 139200 75280
rect 798 74736 139200 75000
rect 880 74456 139200 74736
rect 798 74192 139200 74456
rect 880 73912 139200 74192
rect 798 73648 139200 73912
rect 880 73368 139200 73648
rect 798 73104 139200 73368
rect 880 72824 139200 73104
rect 798 72560 139200 72824
rect 880 72288 139200 72560
rect 880 72280 139120 72288
rect 798 72016 139120 72280
rect 880 72008 139120 72016
rect 880 71736 139200 72008
rect 798 71472 139200 71736
rect 880 71192 139200 71472
rect 798 70928 139200 71192
rect 880 70648 139200 70928
rect 798 70384 139200 70648
rect 880 70104 139200 70384
rect 798 69840 139200 70104
rect 880 69560 139200 69840
rect 798 69296 139200 69560
rect 880 69016 139200 69296
rect 798 68752 139200 69016
rect 880 68472 139200 68752
rect 798 68208 139200 68472
rect 880 67928 139200 68208
rect 798 67664 139200 67928
rect 880 67384 139120 67664
rect 798 67120 139200 67384
rect 880 66840 139200 67120
rect 798 66576 139200 66840
rect 880 66296 139200 66576
rect 798 66032 139200 66296
rect 880 65752 139200 66032
rect 798 65488 139200 65752
rect 880 65208 139200 65488
rect 798 64944 139200 65208
rect 880 64664 139200 64944
rect 798 64400 139200 64664
rect 880 64120 139200 64400
rect 798 63856 139200 64120
rect 880 63576 139200 63856
rect 798 63312 139200 63576
rect 880 63040 139200 63312
rect 880 63032 139120 63040
rect 798 62768 139120 63032
rect 880 62760 139120 62768
rect 880 62488 139200 62760
rect 798 62224 139200 62488
rect 880 61944 139200 62224
rect 798 61680 139200 61944
rect 880 61400 139200 61680
rect 798 61136 139200 61400
rect 880 60856 139200 61136
rect 798 60592 139200 60856
rect 880 60312 139200 60592
rect 798 60048 139200 60312
rect 880 59768 139200 60048
rect 798 59504 139200 59768
rect 880 59224 139200 59504
rect 798 58960 139200 59224
rect 880 58680 139200 58960
rect 798 58416 139200 58680
rect 880 58136 139120 58416
rect 798 57872 139200 58136
rect 880 57592 139200 57872
rect 798 57328 139200 57592
rect 880 57048 139200 57328
rect 798 56784 139200 57048
rect 880 56504 139200 56784
rect 798 56240 139200 56504
rect 880 55960 139200 56240
rect 798 55696 139200 55960
rect 880 55416 139200 55696
rect 798 55152 139200 55416
rect 880 54872 139200 55152
rect 798 54608 139200 54872
rect 880 54328 139200 54608
rect 798 54064 139200 54328
rect 880 53792 139200 54064
rect 880 53784 139120 53792
rect 798 53520 139120 53784
rect 880 53512 139120 53520
rect 880 53240 139200 53512
rect 798 52976 139200 53240
rect 880 52696 139200 52976
rect 798 52432 139200 52696
rect 880 52152 139200 52432
rect 798 51888 139200 52152
rect 880 51608 139200 51888
rect 798 51344 139200 51608
rect 880 51064 139200 51344
rect 798 50800 139200 51064
rect 880 50520 139200 50800
rect 798 50256 139200 50520
rect 880 49976 139200 50256
rect 798 49712 139200 49976
rect 880 49432 139200 49712
rect 798 49168 139200 49432
rect 880 48888 139120 49168
rect 798 48624 139200 48888
rect 880 48344 139200 48624
rect 798 48080 139200 48344
rect 880 47800 139200 48080
rect 798 47536 139200 47800
rect 880 47256 139200 47536
rect 798 46992 139200 47256
rect 880 46712 139200 46992
rect 798 46448 139200 46712
rect 880 46168 139200 46448
rect 798 45904 139200 46168
rect 880 45624 139200 45904
rect 798 45360 139200 45624
rect 880 45080 139200 45360
rect 798 44816 139200 45080
rect 880 44544 139200 44816
rect 880 44536 139120 44544
rect 798 44272 139120 44536
rect 880 44264 139120 44272
rect 880 43992 139200 44264
rect 798 43728 139200 43992
rect 880 43448 139200 43728
rect 798 43184 139200 43448
rect 880 42904 139200 43184
rect 798 42640 139200 42904
rect 880 42360 139200 42640
rect 798 42096 139200 42360
rect 880 41816 139200 42096
rect 798 41552 139200 41816
rect 880 41272 139200 41552
rect 798 41008 139200 41272
rect 880 40728 139200 41008
rect 798 40464 139200 40728
rect 880 40184 139200 40464
rect 798 39920 139200 40184
rect 880 39640 139120 39920
rect 798 39376 139200 39640
rect 880 39096 139200 39376
rect 798 38832 139200 39096
rect 880 38552 139200 38832
rect 798 38288 139200 38552
rect 880 38008 139200 38288
rect 798 37744 139200 38008
rect 880 37464 139200 37744
rect 798 37200 139200 37464
rect 880 36920 139200 37200
rect 798 36656 139200 36920
rect 880 36376 139200 36656
rect 798 36112 139200 36376
rect 880 35832 139200 36112
rect 798 35568 139200 35832
rect 880 35296 139200 35568
rect 880 35288 139120 35296
rect 798 35024 139120 35288
rect 880 35016 139120 35024
rect 880 34744 139200 35016
rect 798 34480 139200 34744
rect 880 34200 139200 34480
rect 798 33936 139200 34200
rect 880 33656 139200 33936
rect 798 33392 139200 33656
rect 880 33112 139200 33392
rect 798 32848 139200 33112
rect 880 32568 139200 32848
rect 798 32304 139200 32568
rect 880 32024 139200 32304
rect 798 31760 139200 32024
rect 880 31480 139200 31760
rect 798 31216 139200 31480
rect 880 30936 139200 31216
rect 798 30672 139200 30936
rect 880 30392 139120 30672
rect 798 30128 139200 30392
rect 880 29848 139200 30128
rect 798 29584 139200 29848
rect 880 29304 139200 29584
rect 798 29040 139200 29304
rect 880 28760 139200 29040
rect 798 28496 139200 28760
rect 880 28216 139200 28496
rect 798 27952 139200 28216
rect 880 27672 139200 27952
rect 798 27408 139200 27672
rect 880 27128 139200 27408
rect 798 26864 139200 27128
rect 880 26584 139200 26864
rect 798 26320 139200 26584
rect 880 26048 139200 26320
rect 880 26040 139120 26048
rect 798 25776 139120 26040
rect 880 25768 139120 25776
rect 880 25496 139200 25768
rect 798 25232 139200 25496
rect 880 24952 139200 25232
rect 798 24688 139200 24952
rect 880 24408 139200 24688
rect 798 24144 139200 24408
rect 880 23864 139200 24144
rect 798 23600 139200 23864
rect 880 23320 139200 23600
rect 798 23056 139200 23320
rect 880 22776 139200 23056
rect 798 22512 139200 22776
rect 880 22232 139200 22512
rect 798 21968 139200 22232
rect 880 21688 139200 21968
rect 798 21424 139200 21688
rect 880 21144 139120 21424
rect 798 20880 139200 21144
rect 880 20600 139200 20880
rect 798 20336 139200 20600
rect 880 20056 139200 20336
rect 798 19792 139200 20056
rect 880 19512 139200 19792
rect 798 19248 139200 19512
rect 880 18968 139200 19248
rect 798 18704 139200 18968
rect 880 18424 139200 18704
rect 798 18160 139200 18424
rect 880 17880 139200 18160
rect 798 17616 139200 17880
rect 880 17336 139200 17616
rect 798 17072 139200 17336
rect 880 16800 139200 17072
rect 880 16792 139120 16800
rect 798 16528 139120 16792
rect 880 16520 139120 16528
rect 880 16248 139200 16520
rect 798 15984 139200 16248
rect 880 15704 139200 15984
rect 798 15440 139200 15704
rect 880 15160 139200 15440
rect 798 14896 139200 15160
rect 880 14616 139200 14896
rect 798 14352 139200 14616
rect 880 14072 139200 14352
rect 798 13808 139200 14072
rect 880 13528 139200 13808
rect 798 13264 139200 13528
rect 880 12984 139200 13264
rect 798 12720 139200 12984
rect 880 12440 139200 12720
rect 798 12176 139200 12440
rect 880 11896 139120 12176
rect 798 11632 139200 11896
rect 880 11352 139200 11632
rect 798 11088 139200 11352
rect 880 10808 139200 11088
rect 798 7552 139200 10808
rect 798 7272 139120 7552
rect 798 2928 139200 7272
rect 798 2648 139120 2928
rect 798 2143 139200 2648
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 4843 7787 8221 129845
<< labels >>
rlabel metal2 s 3146 139200 3202 140000 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal2 s 36542 139200 36598 140000 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal2 s 39578 139200 39634 140000 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal2 s 42614 139200 42670 140000 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal2 s 45650 139200 45706 140000 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal2 s 48686 139200 48742 140000 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal2 s 51722 139200 51778 140000 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal2 s 54758 139200 54814 140000 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal2 s 57794 139200 57850 140000 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal2 s 60830 139200 60886 140000 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal2 s 63866 139200 63922 140000 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal2 s 7194 139200 7250 140000 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal2 s 66902 139200 66958 140000 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal2 s 69938 139200 69994 140000 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal2 s 72974 139200 73030 140000 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal2 s 76010 139200 76066 140000 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal2 s 79046 139200 79102 140000 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal2 s 82082 139200 82138 140000 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal2 s 85118 139200 85174 140000 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal2 s 88154 139200 88210 140000 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal2 s 91190 139200 91246 140000 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal2 s 94226 139200 94282 140000 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal2 s 11242 139200 11298 140000 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal2 s 97262 139200 97318 140000 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal2 s 100298 139200 100354 140000 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal2 s 15290 139200 15346 140000 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal2 s 18326 139200 18382 140000 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal2 s 21362 139200 21418 140000 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal2 s 24398 139200 24454 140000 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal2 s 27434 139200 27490 140000 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal2 s 30470 139200 30526 140000 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal2 s 33506 139200 33562 140000 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal2 s 4158 139200 4214 140000 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal2 s 37554 139200 37610 140000 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal2 s 40590 139200 40646 140000 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal2 s 43626 139200 43682 140000 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal2 s 46662 139200 46718 140000 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal2 s 49698 139200 49754 140000 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal2 s 52734 139200 52790 140000 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal2 s 55770 139200 55826 140000 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal2 s 58806 139200 58862 140000 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal2 s 61842 139200 61898 140000 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal2 s 64878 139200 64934 140000 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal2 s 8206 139200 8262 140000 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal2 s 67914 139200 67970 140000 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal2 s 70950 139200 71006 140000 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal2 s 73986 139200 74042 140000 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal2 s 77022 139200 77078 140000 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal2 s 80058 139200 80114 140000 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal2 s 83094 139200 83150 140000 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal2 s 86130 139200 86186 140000 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal2 s 89166 139200 89222 140000 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal2 s 92202 139200 92258 140000 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal2 s 95238 139200 95294 140000 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal2 s 12254 139200 12310 140000 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal2 s 98274 139200 98330 140000 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal2 s 101310 139200 101366 140000 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal2 s 16302 139200 16358 140000 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal2 s 19338 139200 19394 140000 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal2 s 22374 139200 22430 140000 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal2 s 25410 139200 25466 140000 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal2 s 28446 139200 28502 140000 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal2 s 31482 139200 31538 140000 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal2 s 34518 139200 34574 140000 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal2 s 5170 139200 5226 140000 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal2 s 38566 139200 38622 140000 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal2 s 41602 139200 41658 140000 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal2 s 44638 139200 44694 140000 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal2 s 47674 139200 47730 140000 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal2 s 50710 139200 50766 140000 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal2 s 53746 139200 53802 140000 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal2 s 56782 139200 56838 140000 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal2 s 59818 139200 59874 140000 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal2 s 62854 139200 62910 140000 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal2 s 65890 139200 65946 140000 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal2 s 9218 139200 9274 140000 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal2 s 68926 139200 68982 140000 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal2 s 71962 139200 72018 140000 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal2 s 74998 139200 75054 140000 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal2 s 78034 139200 78090 140000 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal2 s 81070 139200 81126 140000 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal2 s 84106 139200 84162 140000 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal2 s 87142 139200 87198 140000 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal2 s 90178 139200 90234 140000 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal2 s 93214 139200 93270 140000 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal2 s 96250 139200 96306 140000 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal2 s 13266 139200 13322 140000 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal2 s 99286 139200 99342 140000 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal2 s 102322 139200 102378 140000 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal2 s 17314 139200 17370 140000 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal2 s 20350 139200 20406 140000 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal2 s 23386 139200 23442 140000 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal2 s 26422 139200 26478 140000 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal2 s 29458 139200 29514 140000 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal2 s 32494 139200 32550 140000 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal2 s 35530 139200 35586 140000 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal2 s 6182 139200 6238 140000 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal2 s 10230 139200 10286 140000 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal2 s 14278 139200 14334 140000 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal3 s 139200 7352 140000 7472 6 io_oeb[0]
port 100 nsew signal output
rlabel metal3 s 139200 99832 140000 99952 6 io_oeb[10]
port 101 nsew signal output
rlabel metal3 s 139200 109080 140000 109200 6 io_oeb[11]
port 102 nsew signal output
rlabel metal3 s 139200 118328 140000 118448 6 io_oeb[12]
port 103 nsew signal output
rlabel metal3 s 139200 127576 140000 127696 6 io_oeb[13]
port 104 nsew signal output
rlabel metal3 s 139200 136824 140000 136944 6 io_oeb[14]
port 105 nsew signal output
rlabel metal2 s 136730 139200 136786 140000 6 io_oeb[15]
port 106 nsew signal output
rlabel metal2 s 134706 139200 134762 140000 6 io_oeb[16]
port 107 nsew signal output
rlabel metal2 s 132682 139200 132738 140000 6 io_oeb[17]
port 108 nsew signal output
rlabel metal2 s 130658 139200 130714 140000 6 io_oeb[18]
port 109 nsew signal output
rlabel metal2 s 128634 139200 128690 140000 6 io_oeb[19]
port 110 nsew signal output
rlabel metal3 s 139200 16600 140000 16720 6 io_oeb[1]
port 111 nsew signal output
rlabel metal2 s 126610 139200 126666 140000 6 io_oeb[20]
port 112 nsew signal output
rlabel metal2 s 124586 139200 124642 140000 6 io_oeb[21]
port 113 nsew signal output
rlabel metal2 s 122562 139200 122618 140000 6 io_oeb[22]
port 114 nsew signal output
rlabel metal2 s 120538 139200 120594 140000 6 io_oeb[23]
port 115 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 io_oeb[24]
port 116 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 io_oeb[25]
port 117 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 io_oeb[26]
port 118 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 io_oeb[27]
port 119 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 io_oeb[28]
port 120 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 io_oeb[29]
port 121 nsew signal output
rlabel metal3 s 139200 25848 140000 25968 6 io_oeb[2]
port 122 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 io_oeb[30]
port 123 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 io_oeb[31]
port 124 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 io_oeb[32]
port 125 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 io_oeb[33]
port 126 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 io_oeb[34]
port 127 nsew signal output
rlabel metal3 s 0 126760 800 126880 6 io_oeb[35]
port 128 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 io_oeb[36]
port 129 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 io_oeb[37]
port 130 nsew signal output
rlabel metal3 s 139200 35096 140000 35216 6 io_oeb[3]
port 131 nsew signal output
rlabel metal3 s 139200 44344 140000 44464 6 io_oeb[4]
port 132 nsew signal output
rlabel metal3 s 139200 53592 140000 53712 6 io_oeb[5]
port 133 nsew signal output
rlabel metal3 s 139200 62840 140000 62960 6 io_oeb[6]
port 134 nsew signal output
rlabel metal3 s 139200 72088 140000 72208 6 io_oeb[7]
port 135 nsew signal output
rlabel metal3 s 139200 81336 140000 81456 6 io_oeb[8]
port 136 nsew signal output
rlabel metal3 s 139200 90584 140000 90704 6 io_oeb[9]
port 137 nsew signal output
rlabel metal3 s 139200 2728 140000 2848 6 io_out[0]
port 138 nsew signal output
rlabel metal3 s 139200 95208 140000 95328 6 io_out[10]
port 139 nsew signal output
rlabel metal3 s 139200 104456 140000 104576 6 io_out[11]
port 140 nsew signal output
rlabel metal3 s 139200 113704 140000 113824 6 io_out[12]
port 141 nsew signal output
rlabel metal3 s 139200 122952 140000 123072 6 io_out[13]
port 142 nsew signal output
rlabel metal3 s 139200 132200 140000 132320 6 io_out[14]
port 143 nsew signal output
rlabel metal2 s 135718 139200 135774 140000 6 io_out[15]
port 144 nsew signal output
rlabel metal2 s 133694 139200 133750 140000 6 io_out[16]
port 145 nsew signal output
rlabel metal2 s 131670 139200 131726 140000 6 io_out[17]
port 146 nsew signal output
rlabel metal2 s 129646 139200 129702 140000 6 io_out[18]
port 147 nsew signal output
rlabel metal2 s 127622 139200 127678 140000 6 io_out[19]
port 148 nsew signal output
rlabel metal3 s 139200 11976 140000 12096 6 io_out[1]
port 149 nsew signal output
rlabel metal2 s 125598 139200 125654 140000 6 io_out[20]
port 150 nsew signal output
rlabel metal2 s 123574 139200 123630 140000 6 io_out[21]
port 151 nsew signal output
rlabel metal2 s 121550 139200 121606 140000 6 io_out[22]
port 152 nsew signal output
rlabel metal2 s 119526 139200 119582 140000 6 io_out[23]
port 153 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 io_out[24]
port 154 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 io_out[25]
port 155 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 io_out[26]
port 156 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 io_out[27]
port 157 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 io_out[28]
port 158 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 io_out[29]
port 159 nsew signal output
rlabel metal3 s 139200 21224 140000 21344 6 io_out[2]
port 160 nsew signal output
rlabel metal3 s 0 120776 800 120896 6 io_out[30]
port 161 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 io_out[31]
port 162 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 io_out[32]
port 163 nsew signal output
rlabel metal3 s 0 124040 800 124160 6 io_out[33]
port 164 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 io_out[34]
port 165 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 io_out[35]
port 166 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 io_out[36]
port 167 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 io_out[37]
port 168 nsew signal output
rlabel metal3 s 139200 30472 140000 30592 6 io_out[3]
port 169 nsew signal output
rlabel metal3 s 139200 39720 140000 39840 6 io_out[4]
port 170 nsew signal output
rlabel metal3 s 139200 48968 140000 49088 6 io_out[5]
port 171 nsew signal output
rlabel metal3 s 139200 58216 140000 58336 6 io_out[6]
port 172 nsew signal output
rlabel metal3 s 139200 67464 140000 67584 6 io_out[7]
port 173 nsew signal output
rlabel metal3 s 139200 76712 140000 76832 6 io_out[8]
port 174 nsew signal output
rlabel metal3 s 139200 85960 140000 86080 6 io_out[9]
port 175 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 mem0_data_i[0]
port 176 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 mem0_data_i[10]
port 177 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 mem0_data_i[11]
port 178 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 mem0_data_i[12]
port 179 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 mem0_data_i[13]
port 180 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 mem0_data_i[14]
port 181 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 mem0_data_i[15]
port 182 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 mem0_data_i[16]
port 183 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 mem0_data_i[17]
port 184 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 mem0_data_i[18]
port 185 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 mem0_data_i[19]
port 186 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 mem0_data_i[1]
port 187 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 mem0_data_i[20]
port 188 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 mem0_data_i[21]
port 189 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 mem0_data_i[22]
port 190 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 mem0_data_i[23]
port 191 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 mem0_data_i[24]
port 192 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 mem0_data_i[25]
port 193 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 mem0_data_i[26]
port 194 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 mem0_data_i[27]
port 195 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 mem0_data_i[28]
port 196 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 mem0_data_i[29]
port 197 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 mem0_data_i[2]
port 198 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 mem0_data_i[30]
port 199 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 mem0_data_i[31]
port 200 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 mem0_data_i[3]
port 201 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 mem0_data_i[4]
port 202 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 mem0_data_i[5]
port 203 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 mem0_data_i[6]
port 204 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 mem0_data_i[7]
port 205 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 mem0_data_i[8]
port 206 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 mem0_data_i[9]
port 207 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 mem1_data_i[0]
port 208 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 mem1_data_i[10]
port 209 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 mem1_data_i[11]
port 210 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 mem1_data_i[12]
port 211 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 mem1_data_i[13]
port 212 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 mem1_data_i[14]
port 213 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 mem1_data_i[15]
port 214 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 mem1_data_i[16]
port 215 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 mem1_data_i[17]
port 216 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mem1_data_i[18]
port 217 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 mem1_data_i[19]
port 218 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 mem1_data_i[1]
port 219 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 mem1_data_i[20]
port 220 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 mem1_data_i[21]
port 221 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 mem1_data_i[22]
port 222 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 mem1_data_i[23]
port 223 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 mem1_data_i[24]
port 224 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 mem1_data_i[25]
port 225 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 mem1_data_i[26]
port 226 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 mem1_data_i[27]
port 227 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 mem1_data_i[28]
port 228 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 mem1_data_i[29]
port 229 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 mem1_data_i[2]
port 230 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 mem1_data_i[30]
port 231 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 mem1_data_i[31]
port 232 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 mem1_data_i[3]
port 233 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 mem1_data_i[4]
port 234 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 mem1_data_i[5]
port 235 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 mem1_data_i[6]
port 236 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 mem1_data_i[7]
port 237 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 mem1_data_i[8]
port 238 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 mem1_data_i[9]
port 239 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 mem2_data_i[0]
port 240 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 mem2_data_i[10]
port 241 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 mem2_data_i[11]
port 242 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 mem2_data_i[12]
port 243 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 mem2_data_i[13]
port 244 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 mem2_data_i[14]
port 245 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 mem2_data_i[15]
port 246 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 mem2_data_i[16]
port 247 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 mem2_data_i[17]
port 248 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 mem2_data_i[18]
port 249 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 mem2_data_i[19]
port 250 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 mem2_data_i[1]
port 251 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 mem2_data_i[20]
port 252 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 mem2_data_i[21]
port 253 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 mem2_data_i[22]
port 254 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 mem2_data_i[23]
port 255 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 mem2_data_i[24]
port 256 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 mem2_data_i[25]
port 257 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 mem2_data_i[26]
port 258 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 mem2_data_i[27]
port 259 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 mem2_data_i[28]
port 260 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 mem2_data_i[29]
port 261 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 mem2_data_i[2]
port 262 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 mem2_data_i[30]
port 263 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 mem2_data_i[31]
port 264 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 mem2_data_i[3]
port 265 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 mem2_data_i[4]
port 266 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 mem2_data_i[5]
port 267 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 mem2_data_i[6]
port 268 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 mem2_data_i[7]
port 269 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 mem2_data_i[8]
port 270 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 mem2_data_i[9]
port 271 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 mem3_data_i[0]
port 272 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 mem3_data_i[10]
port 273 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mem3_data_i[11]
port 274 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 mem3_data_i[12]
port 275 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 mem3_data_i[13]
port 276 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 mem3_data_i[14]
port 277 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 mem3_data_i[15]
port 278 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 mem3_data_i[16]
port 279 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 mem3_data_i[17]
port 280 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 mem3_data_i[18]
port 281 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 mem3_data_i[19]
port 282 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 mem3_data_i[1]
port 283 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 mem3_data_i[20]
port 284 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 mem3_data_i[21]
port 285 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 mem3_data_i[22]
port 286 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 mem3_data_i[23]
port 287 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 mem3_data_i[24]
port 288 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 mem3_data_i[25]
port 289 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 mem3_data_i[26]
port 290 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 mem3_data_i[27]
port 291 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 mem3_data_i[28]
port 292 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 mem3_data_i[29]
port 293 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 mem3_data_i[2]
port 294 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 mem3_data_i[30]
port 295 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 mem3_data_i[31]
port 296 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 mem3_data_i[3]
port 297 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 mem3_data_i[4]
port 298 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 mem3_data_i[5]
port 299 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 mem3_data_i[6]
port 300 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 mem3_data_i[7]
port 301 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 mem3_data_i[8]
port 302 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 mem3_data_i[9]
port 303 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mem_data_o[0]
port 304 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 mem_data_o[10]
port 305 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 mem_data_o[11]
port 306 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 mem_data_o[12]
port 307 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 mem_data_o[13]
port 308 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 mem_data_o[14]
port 309 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 mem_data_o[15]
port 310 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 mem_data_o[16]
port 311 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 mem_data_o[17]
port 312 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 mem_data_o[18]
port 313 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 mem_data_o[19]
port 314 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 mem_data_o[1]
port 315 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 mem_data_o[20]
port 316 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 mem_data_o[21]
port 317 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 mem_data_o[22]
port 318 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 mem_data_o[23]
port 319 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 mem_data_o[24]
port 320 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 mem_data_o[25]
port 321 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 mem_data_o[26]
port 322 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 mem_data_o[27]
port 323 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 mem_data_o[28]
port 324 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 mem_data_o[29]
port 325 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 mem_data_o[2]
port 326 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 mem_data_o[30]
port 327 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 mem_data_o[31]
port 328 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 mem_data_o[3]
port 329 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 mem_data_o[4]
port 330 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 mem_data_o[5]
port 331 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 mem_data_o[6]
port 332 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 mem_data_o[7]
port 333 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 mem_data_o[8]
port 334 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 mem_data_o[9]
port 335 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 mem_raddr_o[0]
port 336 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 mem_raddr_o[1]
port 337 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 mem_raddr_o[2]
port 338 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 mem_raddr_o[3]
port 339 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 mem_raddr_o[4]
port 340 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 mem_raddr_o[5]
port 341 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 mem_raddr_o[6]
port 342 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 mem_raddr_o[7]
port 343 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 mem_raddr_o[8]
port 344 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 mem_renb_o[0]
port 345 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 mem_renb_o[1]
port 346 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 mem_renb_o[2]
port 347 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 mem_renb_o[3]
port 348 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 mem_waddr_o[0]
port 349 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 mem_waddr_o[1]
port 350 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 mem_waddr_o[2]
port 351 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 mem_waddr_o[3]
port 352 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 mem_waddr_o[4]
port 353 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 mem_waddr_o[5]
port 354 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 mem_waddr_o[6]
port 355 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 mem_waddr_o[7]
port 356 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 mem_waddr_o[8]
port 357 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 mem_wenb_o[0]
port 358 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 mem_wenb_o[1]
port 359 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 mem_wenb_o[2]
port 360 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 mem_wenb_o[3]
port 361 nsew signal output
rlabel metal2 s 103334 139200 103390 140000 6 oversample_o[0]
port 362 nsew signal output
rlabel metal2 s 104346 139200 104402 140000 6 oversample_o[1]
port 363 nsew signal output
rlabel metal2 s 105358 139200 105414 140000 6 oversample_o[2]
port 364 nsew signal output
rlabel metal2 s 106370 139200 106426 140000 6 oversample_o[3]
port 365 nsew signal output
rlabel metal2 s 107382 139200 107438 140000 6 oversample_o[4]
port 366 nsew signal output
rlabel metal2 s 108394 139200 108450 140000 6 oversample_o[5]
port 367 nsew signal output
rlabel metal2 s 109406 139200 109462 140000 6 oversample_o[6]
port 368 nsew signal output
rlabel metal2 s 110418 139200 110474 140000 6 oversample_o[7]
port 369 nsew signal output
rlabel metal2 s 111430 139200 111486 140000 6 oversample_o[8]
port 370 nsew signal output
rlabel metal2 s 112442 139200 112498 140000 6 oversample_o[9]
port 371 nsew signal output
rlabel metal2 s 116490 139200 116546 140000 6 sinc3_en_o[0]
port 372 nsew signal output
rlabel metal2 s 117502 139200 117558 140000 6 sinc3_en_o[1]
port 373 nsew signal output
rlabel metal2 s 118514 139200 118570 140000 6 sinc3_en_o[2]
port 374 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 375 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 375 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 375 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 375 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 375 nsew power bidirectional
rlabel metal2 s 113454 139200 113510 140000 6 vco_enb_o[0]
port 376 nsew signal output
rlabel metal2 s 114466 139200 114522 140000 6 vco_enb_o[1]
port 377 nsew signal output
rlabel metal2 s 115478 139200 115534 140000 6 vco_enb_o[2]
port 378 nsew signal output
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 379 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 379 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 379 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 379 nsew ground bidirectional
rlabel metal2 s 2318 0 2374 800 6 wb_clk_i
port 380 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wb_rst_i
port 381 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_ack_o
port 382 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[0]
port 383 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_adr_i[10]
port 384 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[11]
port 385 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_adr_i[12]
port 386 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_adr_i[13]
port 387 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[14]
port 388 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[15]
port 389 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_adr_i[16]
port 390 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 wbs_adr_i[17]
port 391 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_adr_i[18]
port 392 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 wbs_adr_i[19]
port 393 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[1]
port 394 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_adr_i[20]
port 395 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 wbs_adr_i[21]
port 396 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_adr_i[22]
port 397 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 wbs_adr_i[23]
port 398 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 wbs_adr_i[24]
port 399 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 wbs_adr_i[25]
port 400 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 wbs_adr_i[26]
port 401 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 wbs_adr_i[27]
port 402 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 wbs_adr_i[28]
port 403 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 wbs_adr_i[29]
port 404 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[2]
port 405 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 wbs_adr_i[30]
port 406 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 wbs_adr_i[31]
port 407 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[3]
port 408 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[4]
port 409 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[5]
port 410 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_adr_i[6]
port 411 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_adr_i[7]
port 412 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[8]
port 413 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_adr_i[9]
port 414 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_cyc_i
port 415 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[0]
port 416 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[10]
port 417 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_dat_i[11]
port 418 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[12]
port 419 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_i[13]
port 420 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_dat_i[14]
port 421 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_i[15]
port 422 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_i[16]
port 423 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_dat_i[17]
port 424 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_i[18]
port 425 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[19]
port 426 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[1]
port 427 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_dat_i[20]
port 428 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_i[21]
port 429 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_i[22]
port 430 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 wbs_dat_i[23]
port 431 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 wbs_dat_i[24]
port 432 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_i[25]
port 433 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 wbs_dat_i[26]
port 434 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 wbs_dat_i[27]
port 435 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 wbs_dat_i[28]
port 436 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 wbs_dat_i[29]
port 437 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[2]
port 438 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 wbs_dat_i[30]
port 439 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 wbs_dat_i[31]
port 440 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[3]
port 441 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[4]
port 442 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_i[5]
port 443 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[6]
port 444 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_i[7]
port 445 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[8]
port 446 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_i[9]
port 447 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[0]
port 448 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_o[10]
port 449 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_o[11]
port 450 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[12]
port 451 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 wbs_dat_o[13]
port 452 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_o[14]
port 453 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 wbs_dat_o[15]
port 454 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[16]
port 455 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 wbs_dat_o[17]
port 456 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 wbs_dat_o[18]
port 457 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 wbs_dat_o[19]
port 458 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[1]
port 459 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_o[20]
port 460 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 wbs_dat_o[21]
port 461 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_o[22]
port 462 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 wbs_dat_o[23]
port 463 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_o[24]
port 464 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_o[25]
port 465 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 wbs_dat_o[26]
port 466 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 wbs_dat_o[27]
port 467 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 wbs_dat_o[28]
port 468 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 wbs_dat_o[29]
port 469 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[2]
port 470 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 wbs_dat_o[30]
port 471 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 wbs_dat_o[31]
port 472 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[3]
port 473 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[4]
port 474 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[5]
port 475 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[6]
port 476 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[7]
port 477 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_o[8]
port 478 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 wbs_dat_o[9]
port 479 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_sel_i[0]
port 480 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_sel_i[1]
port 481 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_sel_i[2]
port 482 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_sel_i[3]
port 483 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_stb_i
port 484 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_we_i
port 485 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 wmask_o[0]
port 486 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 wmask_o[1]
port 487 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 wmask_o[2]
port 488 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 wmask_o[3]
port 489 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8845790
string GDS_FILE /home/cass/work/caravel_vco_adc/openlane/vco_adc_wrapper/runs/23_09_19_16_06/results/signoff/vco_adc_wrapper.magic.gds
string GDS_START 486552
<< end >>

